magic
tech scmos
timestamp 1700521624
<< metal1 >>
rect 127 344 487 348
rect 577 340 606 343
rect 591 325 597 337
rect 96 135 103 142
rect 577 99 606 102
rect 591 83 597 95
rect 76 13 83 20
rect 523 11 530 20
rect -290 -84 -279 -48
rect 157 -55 165 -49
rect 108 -111 116 -92
rect 555 -111 563 -92
rect 578 -139 607 -136
rect 591 -154 597 -142
rect 577 -384 606 -381
rect 591 -401 597 -389
rect 76 -445 83 -435
rect 524 -443 531 -428
rect 398 -548 405 -533
rect 537 -553 558 -547
<< m2contact >>
rect 601 170 609 176
rect 543 110 550 121
rect 938 7 950 17
rect 601 -72 609 -65
rect 564 -88 571 -82
rect 938 -224 950 -214
rect 601 -313 609 -303
rect 96 -327 103 -320
rect 941 -469 950 -458
rect 564 -543 572 -533
rect 601 -551 610 -542
<< metal2 >>
rect -277 318 -271 335
rect 170 318 176 335
rect 547 164 556 198
rect 601 164 609 170
rect 547 157 609 164
rect 157 149 166 156
rect -28 -87 -18 -66
rect 185 -74 191 -57
rect 938 -71 950 7
rect 601 -82 609 -72
rect -28 -97 144 -87
rect 571 -88 609 -82
rect 802 -84 950 -71
rect -277 -137 -271 -120
rect 134 -320 144 -97
rect 802 -115 815 -84
rect 171 -137 177 -120
rect 455 -127 815 -115
rect 938 -214 950 -120
rect 548 -307 557 -258
rect 548 -313 601 -307
rect 103 -327 144 -320
rect 461 -331 496 -320
rect 573 -345 950 -333
rect 941 -458 950 -345
rect 572 -542 610 -533
rect 572 -543 601 -542
<< m3contact >>
rect 382 -74 390 -66
rect 456 -331 461 -320
rect 496 -331 501 -320
rect 558 -345 573 -333
<< m123contact >>
rect 939 251 950 258
rect 587 185 597 194
rect 591 -14 597 -8
rect -58 -55 -48 -47
rect 157 -64 165 -55
rect -290 -93 -279 -84
rect -290 -323 -279 -315
rect 591 -252 597 -246
rect 157 -322 165 -314
rect 544 -345 551 -335
rect 591 -497 597 -491
rect -28 -529 -18 -521
<< metal3 >>
rect 581 -8 587 194
rect 939 149 950 251
rect 624 137 950 149
rect 581 -14 591 -8
rect -58 -64 157 -55
rect -290 -315 -279 -93
rect 157 -314 165 -64
rect 382 -99 390 -74
rect 581 -99 587 -14
rect 382 -107 587 -99
rect 582 -246 588 -107
rect 582 -252 591 -246
rect 391 -331 456 -320
rect 501 -331 573 -320
rect 558 -333 573 -331
rect 147 -345 450 -335
rect 514 -345 544 -335
rect -28 -530 -18 -529
rect 147 -530 158 -345
rect 582 -491 588 -252
rect 582 -497 591 -491
rect -28 -540 158 -530
<< m234contact >>
rect -119 334 -102 348
rect 157 137 166 149
rect 543 99 550 110
rect -178 -115 -161 -97
rect 938 -120 950 -104
rect 400 -529 408 -521
<< m4contact >>
rect 604 137 624 149
rect 383 -331 391 -320
rect 450 -345 456 -335
rect 507 -345 514 -335
<< metal4 >>
rect -102 334 155 343
rect 144 153 155 334
rect 144 131 153 153
rect 166 137 604 149
rect 144 -38 155 131
rect -178 -78 -161 -77
rect -178 -97 376 -78
rect 359 -104 376 -97
rect 144 -320 155 -115
rect 543 -284 550 99
rect 628 -120 938 -104
rect 400 -292 550 -284
rect 144 -331 383 -320
rect 400 -521 408 -292
rect 456 -345 507 -335
<< m5contact >>
rect 144 -47 155 -38
rect 144 -115 155 -106
rect 359 -121 376 -104
rect 610 -120 628 -104
<< metal5 >>
rect 144 -106 155 -47
rect 376 -120 610 -104
use Full_Adder_t3  Full_Adder_t3_3
timestamp 1699877225
transform 1 0 171 0 1 -321
box -13 -232 411 214
use Full_Adder_t3  Full_Adder_t3_2
timestamp 1699877225
transform 1 0 -277 0 1 -321
box -13 -232 411 214
use Full_Adder_t3  Full_Adder_t3_1
timestamp 1699877225
transform 1 0 170 0 1 134
box -13 -232 411 214
use Full_Adder_t3  Full_Adder_t3_0
timestamp 1699877225
transform 1 0 -277 0 1 134
box -13 -232 411 214
use XOR  XOR_0
timestamp 1699269911
transform 1 0 735 0 1 259
box -144 -89 215 89
use XOR  XOR_2
timestamp 1699269911
transform 1 0 735 0 1 -465
box -144 -89 215 89
use XOR  XOR_3
timestamp 1699269911
transform 1 0 735 0 1 -220
box -144 -89 215 89
use XOR  XOR_1
timestamp 1699269911
transform 1 0 735 0 1 18
box -144 -89 215 89
<< end >>
