module Or_G(Y, A, B);
    input A, B;
    output Y;
    assign Y = A|B;
endmodule