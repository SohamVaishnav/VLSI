module Not_G(Y, A);
    input A;
    output Y;
    assign Y = ~A;
endmodule