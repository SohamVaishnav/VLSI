magic
tech scmos
timestamp 1699636190
<< end >>
