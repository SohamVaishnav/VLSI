.title Ring Oscillator

.include TSMC_180nm.txt
.include NOT.sub
.global gnd 

VDD vdd 0 dc 1.8

X1 in w1 vdd gnd NOT 
X2 w1 w2 vdd gnd NOT
X3 w2 in vdd gnd NOT

.ic v(in) = 0

.control 
run
tran 10u 10n
plot v(w2)
.endc 

.end