magic
tech scmos
timestamp 1700515795
<< metal1 >>
rect 135 17 139 22
rect 135 -50 139 -45
rect 135 -117 139 -112
rect 135 -184 139 -179
<< m2contact >>
rect 67 57 76 64
rect -5 42 4 49
rect 104 0 113 7
rect 61 -7 70 0
rect -5 -23 4 -16
rect 104 -67 113 -60
rect 61 -74 70 -67
rect -5 -90 4 -83
rect 104 -134 113 -127
rect 61 -141 70 -134
rect -5 -157 4 -150
rect 104 -201 113 -194
<< metal2 >>
rect 61 57 67 64
rect -5 -16 4 42
rect -5 -83 4 -23
rect -5 -150 4 -90
rect 61 0 70 57
rect 61 -67 70 -7
rect 61 -134 70 -74
rect 104 -60 113 0
rect 104 -127 113 -67
rect 104 -194 113 -134
use 3_input_AND  3_input_AND_3
timestamp 1700132798
transform 1 0 49 0 1 -162
box -49 -39 90 25
use 3_input_AND  3_input_AND_2
timestamp 1700132798
transform 1 0 49 0 1 -95
box -49 -39 90 25
use 3_input_AND  3_input_AND_1
timestamp 1700132798
transform 1 0 49 0 1 -28
box -49 -39 90 25
use 3_input_AND  3_input_AND_0
timestamp 1700132798
transform 1 0 49 0 1 39
box -49 -39 90 25
<< labels >>
flabel metal1 135 17 139 22 0 FreeSans 9 0 0 0 C0
flabel metal1 135 -50 139 -45 0 FreeSans 9 0 0 0 C1
flabel metal1 135 -117 139 -112 0 FreeSans 9 0 0 0 C2
flabel metal1 135 -184 139 -179 0 FreeSans 9 0 0 0 C3
<< end >>
