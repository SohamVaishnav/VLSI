magic
tech scmos
timestamp 1698776833
<< nwell >>
rect -42 -2 -12 34
rect -1 -2 29 34
rect 40 -2 70 34
<< ntransistor >>
rect -35 -21 -20 -16
rect 6 -21 21 -16
rect 47 -21 62 -16
<< ptransistor >>
rect -35 14 -20 19
rect 6 14 21 19
rect 47 14 62 19
<< ndiffusion >>
rect -35 -16 -20 -15
rect 6 -16 21 -15
rect 47 -16 62 -15
rect -35 -22 -20 -21
rect 6 -22 21 -21
rect 47 -22 62 -21
<< pdiffusion >>
rect -35 19 -20 21
rect 6 19 21 21
rect 47 19 62 21
rect -35 12 -20 14
rect 6 12 21 14
rect 47 12 62 14
<< ndcontact >>
rect -35 -15 -20 -9
rect 6 -15 21 -9
rect 47 -15 62 -9
rect -35 -28 -20 -22
rect 6 -28 21 -22
rect 47 -28 62 -22
<< pdcontact >>
rect -35 21 -20 28
rect 6 21 21 28
rect 47 21 62 28
rect -35 5 -20 12
rect 6 5 21 12
rect 47 5 62 12
<< polysilicon >>
rect -42 14 -35 19
rect -20 14 -12 19
rect -1 14 6 19
rect 21 14 29 19
rect 40 14 47 19
rect 62 14 70 19
rect -42 -16 -38 14
rect -1 -16 3 14
rect 35 -16 40 14
rect -38 -21 -35 -16
rect -20 -21 -13 -16
rect 3 -21 6 -16
rect 21 -21 28 -16
rect 35 -21 47 -16
rect 62 -21 69 -16
<< polycontact >>
rect 35 14 40 19
rect -42 -21 -38 -16
rect -1 -21 3 -16
<< metal1 >>
rect -29 37 56 40
rect -47 34 -26 37
rect -29 28 -26 34
rect 12 31 40 34
rect 12 28 15 31
rect 35 19 40 31
rect 53 28 56 37
rect 30 14 35 19
rect -29 1 -26 5
rect 12 1 15 5
rect -29 -2 15 1
rect 30 -6 34 14
rect -29 -9 34 -6
rect 53 1 56 5
rect 53 -2 71 1
rect 53 -9 56 -2
rect -47 -21 -42 -16
rect -6 -21 -1 -16
rect -29 -31 69 -28
<< end >>
