magic
tech scmos
timestamp 1700494881
<< polysilicon >>
rect 384 -383 388 -353
<< metal1 >>
rect -53 158 -49 163
rect -72 155 -71 158
rect -66 155 -49 158
rect 328 160 375 163
rect 328 119 335 160
rect 567 158 637 168
rect 648 165 871 168
rect 648 158 826 165
rect 814 96 826 158
rect 884 126 889 139
rect 871 123 889 126
rect 884 119 889 123
rect -39 82 -34 87
rect -72 79 -34 82
rect 329 -4 335 46
rect 873 39 889 42
rect 329 -7 387 -4
rect 328 -23 371 -20
rect 328 -64 335 -23
rect 738 -31 745 -20
rect 874 -61 888 -58
rect 329 -187 335 -137
rect 724 -163 730 -137
rect 329 -190 390 -187
rect 822 -197 826 -124
rect -48 -201 -29 -197
rect 152 -201 238 -197
rect 233 -216 238 -201
rect 486 -201 572 -197
rect 722 -201 826 -197
rect 486 -216 490 -201
rect 208 -247 242 -243
rect 800 -247 818 -240
rect 162 -277 169 -260
rect 237 -272 242 -247
rect -45 -288 -32 -278
rect 2 -284 15 -278
rect 43 -284 52 -278
rect 228 -284 288 -280
rect 586 -286 598 -277
rect 638 -284 653 -278
rect 750 -287 756 -260
rect 750 -292 801 -287
rect 149 -301 249 -297
rect 482 -301 609 -297
rect 166 -331 170 -316
rect -22 -365 1 -355
rect 68 -370 72 -355
rect 157 -377 206 -373
rect 220 -377 229 -301
rect 237 -357 242 -339
rect 551 -360 590 -355
rect 619 -359 626 -346
rect 722 -373 726 -357
rect 776 -373 782 -292
rect 326 -377 453 -373
rect 575 -377 606 -373
rect 157 -388 162 -377
rect 601 -388 606 -377
rect 722 -379 782 -373
rect -22 -404 27 -394
rect 158 -413 173 -407
rect 732 -415 738 -407
rect 132 -457 140 -444
rect 425 -443 437 -436
rect 575 -440 586 -415
rect 749 -444 757 -379
rect 684 -453 690 -445
rect 726 -448 757 -444
rect 257 -457 261 -454
rect 567 -457 690 -453
rect 132 -461 263 -457
<< m2contact >>
rect -71 153 -66 158
rect 637 158 648 168
rect 875 163 880 168
rect 884 113 889 119
rect 850 89 855 95
rect -96 77 -91 82
rect 329 77 335 83
rect 724 77 730 82
rect 875 78 880 84
rect -71 69 -66 74
rect 737 57 745 64
rect 247 42 258 49
rect -96 -7 -91 -2
rect 889 37 895 42
rect 850 5 855 11
rect -71 -31 -66 -26
rect 875 -21 880 -16
rect 637 -69 648 -60
rect 888 -65 895 -58
rect 738 -75 745 -69
rect 759 -99 764 -94
rect 850 -95 855 -89
rect -96 -107 -91 -102
rect 329 -106 335 -100
rect 724 -106 730 -101
rect -71 -113 -66 -108
rect 875 -110 880 -105
rect 767 -135 773 -130
rect -96 -189 -91 -184
rect 188 -190 195 -184
rect 724 -168 730 -163
rect 873 -150 880 -144
rect 850 -184 855 -179
rect -54 -204 -48 -197
rect 196 -256 201 -250
rect 787 -256 792 -250
rect 15 -284 23 -278
rect 92 -284 97 -278
rect 135 -284 140 -278
rect 162 -284 169 -277
rect 218 -284 228 -277
rect 653 -284 660 -278
rect 683 -284 688 -278
rect 726 -284 731 -278
rect 801 -292 808 -286
rect -7 -304 -1 -297
rect 166 -316 171 -309
rect 28 -359 33 -353
rect 102 -360 107 -355
rect 68 -377 74 -370
rect 127 -371 133 -363
rect 237 -339 248 -329
rect 755 -332 764 -325
rect 293 -361 300 -353
rect 656 -360 661 -355
rect 691 -360 696 -355
rect 269 -369 276 -362
rect 155 -448 163 -442
<< pm12contact >>
rect 442 -358 450 -351
rect 384 -389 391 -383
<< metal2 >>
rect -96 -2 -91 77
rect -96 -102 -91 -7
rect -96 -184 -91 -107
rect -71 74 -66 153
rect -71 -26 -66 69
rect -71 -108 -66 -31
rect 247 -184 258 42
rect 329 40 335 77
rect 347 53 477 60
rect 292 32 335 40
rect 292 23 302 32
rect 292 -119 302 15
rect 195 -190 258 -184
rect 266 -129 302 -119
rect 329 -100 335 -20
rect 637 -60 648 158
rect 724 64 730 77
rect 724 57 737 64
rect 724 41 730 57
rect 696 34 730 41
rect 850 11 855 89
rect -54 -297 -48 -204
rect 15 -278 23 -190
rect 218 -250 228 -190
rect 266 -194 276 -129
rect 329 -142 335 -106
rect 301 -150 335 -142
rect 724 -75 738 -69
rect 724 -101 730 -75
rect 850 -89 855 5
rect 764 -99 773 -94
rect 724 -143 730 -106
rect 653 -149 730 -143
rect 767 -130 773 -99
rect 653 -235 660 -149
rect 767 -163 773 -135
rect 730 -168 773 -163
rect 767 -179 773 -168
rect 850 -179 855 -95
rect 875 84 880 163
rect 875 -16 880 78
rect 889 32 895 37
rect 875 -105 880 -21
rect 767 -184 850 -179
rect 298 -244 660 -235
rect 201 -256 228 -250
rect 218 -277 228 -256
rect 117 -284 135 -278
rect 169 -284 218 -277
rect -54 -304 -7 -297
rect 15 -353 23 -284
rect 171 -316 206 -309
rect 15 -359 28 -353
rect 219 -362 228 -284
rect 653 -278 660 -244
rect 792 -256 808 -250
rect 688 -284 693 -278
rect 801 -286 808 -256
rect 248 -339 359 -329
rect 764 -332 810 -325
rect 317 -353 408 -346
rect 450 -358 463 -351
rect 127 -373 133 -371
rect 219 -369 269 -362
rect 219 -373 228 -369
rect 127 -379 228 -373
rect 155 -442 163 -379
rect 293 -396 300 -361
rect 453 -368 463 -358
rect 453 -378 645 -368
rect 391 -389 422 -383
rect 293 -402 394 -396
rect 385 -424 394 -402
rect 412 -425 422 -389
rect 801 -425 810 -332
rect 873 -352 880 -150
rect 888 -370 895 -65
rect 412 -434 810 -425
<< m3contact >>
rect 15 -190 23 -182
rect 477 53 485 60
rect 292 15 302 23
rect 329 -20 335 -13
rect 292 -150 301 -142
rect 266 -204 276 -194
rect 290 -244 298 -235
rect 206 -316 213 -309
rect 359 -339 369 -329
rect 310 -353 317 -346
rect 408 -353 415 -346
rect 645 -378 655 -368
rect 385 -435 394 -424
<< m123contact >>
rect -109 113 -104 118
rect -109 29 -104 34
rect -109 -71 -104 -66
rect -109 -155 -104 -150
rect -54 143 -48 148
rect 341 142 347 149
rect -54 47 -48 53
rect -54 -41 -48 -35
rect -54 -136 -48 -130
rect 341 -42 347 -35
rect 837 122 845 129
rect 837 38 845 45
rect 737 14 745 23
rect 738 -20 745 -13
rect 837 -62 845 -55
rect 341 -178 349 -171
rect 837 -153 845 -145
rect 293 -275 300 -268
rect 351 -273 358 -266
rect 408 -276 415 -268
rect -32 -288 -22 -278
rect 34 -284 43 -277
rect -32 -365 -22 -355
rect 541 -292 551 -278
rect 578 -286 586 -277
rect 818 -247 827 -240
rect 619 -346 626 -339
rect -32 -404 -22 -394
rect 541 -360 551 -351
rect 173 -413 180 -407
rect 329 -420 336 -413
rect 592 -404 601 -395
rect 738 -415 746 -407
rect 575 -449 586 -440
<< metal3 >>
rect -109 143 -54 148
rect -109 118 -104 143
rect 347 142 393 149
rect 386 129 393 142
rect 386 122 693 129
rect 700 122 837 129
rect -109 47 -54 53
rect -109 34 -104 47
rect 477 45 485 53
rect 477 38 837 45
rect 302 15 737 23
rect 335 -20 738 -13
rect -109 -41 -54 -35
rect -109 -66 -104 -41
rect 347 -42 379 -35
rect 372 -55 379 -42
rect 372 -62 608 -55
rect 620 -62 837 -55
rect -109 -136 -54 -130
rect -109 -150 -104 -136
rect 83 -150 292 -142
rect 83 -182 91 -150
rect 837 -171 845 -153
rect 179 -178 341 -171
rect 349 -178 845 -171
rect 23 -190 585 -182
rect -32 -204 266 -194
rect 276 -204 491 -194
rect -32 -278 -22 -204
rect 34 -244 290 -235
rect 34 -277 43 -244
rect -32 -355 -22 -288
rect 293 -309 300 -275
rect 213 -316 300 -309
rect 329 -273 351 -266
rect 173 -353 310 -346
rect -32 -394 -22 -365
rect 173 -407 180 -353
rect 329 -413 336 -273
rect 359 -447 369 -339
rect 408 -346 415 -276
rect 481 -284 491 -204
rect 578 -277 585 -190
rect 481 -292 541 -284
rect 541 -351 551 -292
rect 578 -339 585 -286
rect 578 -346 619 -339
rect 541 -375 551 -360
rect 818 -368 827 -247
rect 582 -375 590 -374
rect 541 -383 590 -375
rect 655 -378 827 -368
rect 582 -395 590 -383
rect 582 -404 592 -395
rect 738 -424 746 -415
rect 394 -435 746 -424
rect 359 -449 575 -447
rect 359 -458 586 -449
<< m234contact >>
rect 889 113 895 119
rect 341 53 347 60
rect 889 27 895 32
rect 82 -284 92 -278
rect 106 -284 117 -278
rect 97 -360 102 -355
rect 74 -377 81 -370
rect 693 -284 700 -277
rect 731 -284 738 -278
rect 650 -360 656 -355
rect 686 -360 691 -355
rect 873 -359 880 -352
rect 888 -377 895 -370
<< m4contact >>
rect 693 122 700 129
rect 608 -62 620 -55
rect 171 -178 179 -171
<< metal4 >>
rect 82 151 895 158
rect 82 -278 92 151
rect 106 53 341 60
rect 106 -278 117 53
rect 171 -355 179 -178
rect 608 -284 620 -62
rect 693 -277 700 122
rect 889 119 895 151
rect 889 -278 895 27
rect 738 -284 895 -278
rect 608 -292 656 -284
rect 102 -360 179 -355
rect 650 -355 656 -292
rect 686 -355 873 -352
rect 691 -359 873 -355
rect 81 -377 888 -370
use 3_input_AND  3_input_AND_0
timestamp 1700132798
transform 1 0 72 0 1 -409
box -49 -39 90 25
use AND_2  AND_2_0
timestamp 1698776759
transform 1 0 190 0 1 -420
box -8 -37 143 47
use 4_input_OR  4_input_OR_1
timestamp 1700131117
transform 1 0 239 0 1 -333
box -6 -36 278 37
use 4_input_OR  4_input_OR_0
timestamp 1700131117
transform 1 0 239 0 1 -248
box -6 -36 278 37
use 5_input_AND  5_input_AND_0
timestamp 1699638001
transform 1 0 -41 0 1 -239
box -12 -45 256 42
use XNOR  XNOR_1
timestamp 1699700809
transform 1 0 237 0 1 -160
box -291 -33 98 145
use 4_input_AND  4_input_AND_0
timestamp 1700132235
transform 1 0 61 0 1 -314
box -64 -53 109 17
use 3_input_AND  3_input_AND_1
timestamp 1700132798
transform 1 0 646 0 1 -409
box -49 -39 90 25
use AND_2  AND_2_1
timestamp 1698776759
transform 1 0 438 0 1 -420
box -8 -37 143 47
use 5_input_AND  5_input_AND_1
timestamp 1699638001
transform 1 0 550 0 1 -239
box -12 -45 256 42
use XNOR  XNOR_3
timestamp 1699700809
transform 1 0 632 0 1 -160
box -291 -33 98 145
use 4_input_AND  4_input_AND_1
timestamp 1700132235
transform 1 0 650 0 1 -314
box -64 -53 109 17
use XNOR  XNOR_0
timestamp 1699700809
transform 1 0 237 0 1 23
box -291 -33 98 145
use XNOR  XNOR_2
timestamp 1699700809
transform 1 0 632 0 1 23
box -291 -33 98 145
use 5_input_AND  5_input_AND_2
timestamp 1699638001
transform 0 1 784 -1 0 107
box -12 -45 256 42
use CMOS_in  CMOS_in_7
timestamp 1699269643
transform 1 0 850 0 1 -144
box -13 -40 30 39
use CMOS_in  CMOS_in_6
timestamp 1699269643
transform 1 0 850 0 1 -55
box -13 -40 30 39
use CMOS_in  CMOS_in_5
timestamp 1699269643
transform 1 0 850 0 1 45
box -13 -40 30 39
use CMOS_in  CMOS_in_4
timestamp 1699269643
transform 1 0 850 0 1 129
box -13 -40 30 39
use CMOS_in  CMOS_in_3
timestamp 1699269643
transform 1 0 -96 0 1 -149
box -13 -40 30 39
use CMOS_in  CMOS_in_2
timestamp 1699269643
transform 1 0 -96 0 1 -65
box -13 -40 30 39
use CMOS_in  CMOS_in_1
timestamp 1699269643
transform 1 0 -96 0 1 35
box -13 -40 30 39
use CMOS_in  CMOS_in_0
timestamp 1699269643
transform 1 0 -96 0 1 119
box -13 -40 30 39
<< end >>
