.title Majority Func

.include TSMC_180nm.txt 
.include 4_1_MUX.sub
.global gnd

VA A 0 PULSE(0 1.8 0 100p 100p 20n 40n)
VB B 0 PULSE(0 1.8 0 100p 100p 20n 40n)
VC C 0 PULSE(0 1.8 0 100p 100p 20n 40n)

VDD vdd gnd dc 1.8

X1 A B 0 C C vdd Fn vdd gnd 4_1_MUX

CL Fn 0 2fF

.tran 10u 100n
* .measure tran trise
* + TRIG v(A) VAL = 0.9 RISE =1
* + TARG v(Fn) VAL = 0.9 RISE =1 

* .measure tran tfall
* + TRIG v(A) VAL = 0.9 FALL =1 
* + TARG v(Fn) VAL = 0.9 FALL =1

* .measure tran tpd PARAM = '(trise + tfall)/2' GOAL = 0

* .measure tran triseB
* + TRIG v(B) VAL = 0.9 RISE =1
* + TARG v(Fn) VAL = 0.9 RISE =1 

* .measure tran tfallB
* + TRIG v(B) VAL = 0.9 FALL =1 
* + TARG v(Fn) VAL = 0.9 FALL =1

* .measure tran tpd PARAM = '(triseB + tfallB)/2' GOAL = 0

* .measure tran triseC
* + TRIG v(C) VAL = 0.9 RISE =1
* + TARG v(Fn) VAL = 0.9 RISE =1 

* .measure tran tfallC
* + TRIG v(C) VAL = 0.9 FALL =1 
* + TARG v(Fn) VAL = 0.9 FALL =1

* .measure tran tpd PARAM = '(triseC + tfallC)/2' GOAL = 0

.control 
run 
plot v(Fn) v(A)+2 v(B)+4 v(C)+6
quit
.endc
.end