.title 4 Bit ALU
.include TSMC_180nm.txt
.include NOT.sub
.include NAND.sub
.include NOR.sub
.include AND.sub
.include OR.sub

VinSel0 sel0 0 PULSE(0 3.3 0 100p 100p 10u 20u)
VinSel1 sel1 0 PULSE(0 3.3 0 100p 100p 20u 40u)

*let A be 1010 and B be 1100
VinA inA 0 PULSE(0 3.3 0 100p 100p 10u 20u) 
VinB inB 0 PULSE(0 3.3 0 100p 100p 20u 40u)

VDD vdd 0 3.3

*Decoder
X1 sel0 s0 vdd 0 NOT
X2 sel1 s1 vdd 0 NOT
X3 s0 s1 y1 vdd 0 AND
X4 s0 sel1 y2 vdd 0 AND
X5 sel0 s1 y3 vdd 0 AND
X6 sel0 sel1 y4 vdd 0 AND

*4 bit ANDer
X7 inA inB ANDed vdd 0 AND

.control 
run
tran 10u 40u
plot v(sel0) v(sel1)
plot v(y1) v(y2)+2 v(y3)+4 v(y4)+8
plot v(ANDed)
hardcopy image.ps v(y1) v(y2)+2 v(y3)+4 v(y4)+8
hardcopy image.ps v(ANDed)
.endc

.end