magic
tech scmos
timestamp 1698930095
<< polysilicon >>
rect 531 439 752 450
rect 163 434 167 437
rect 163 416 167 430
rect 743 414 752 439
rect 1082 434 1300 451
rect 1633 434 1841 447
rect 742 407 752 414
rect 1290 407 1300 434
rect 1830 414 1841 434
<< polycontact >>
rect 163 437 167 441
rect 515 439 531 450
rect 163 430 167 434
rect 163 409 167 416
rect 1071 434 1082 451
rect 1619 434 1633 447
rect 730 407 742 414
rect 1279 407 1290 414
rect 1830 407 1841 414
<< metal1 >>
rect 33 632 284 640
rect 582 632 829 640
rect 33 544 45 632
rect 55 590 64 608
rect 165 602 175 610
rect 582 555 593 632
rect 1126 628 1378 636
rect 600 590 609 608
rect 32 540 83 544
rect 33 425 45 540
rect 55 434 61 499
rect 400 459 405 550
rect 234 453 405 459
rect 434 544 593 555
rect 1126 554 1136 628
rect 1676 627 1925 635
rect 1149 586 1158 603
rect 1676 566 1685 627
rect 1696 585 1705 610
rect 434 542 633 544
rect 234 449 244 453
rect 163 441 167 445
rect 55 430 163 434
rect 167 430 193 434
rect 182 429 193 430
rect 0 408 7 425
rect 17 419 114 425
rect 434 419 438 542
rect 582 540 633 542
rect 170 409 183 416
rect 384 408 403 415
rect 117 -19 124 60
rect 195 -8 206 39
rect 515 -8 531 439
rect 582 423 593 540
rect 945 462 950 550
rect 783 455 950 462
rect 983 542 1136 554
rect 1531 553 1685 566
rect 783 447 790 455
rect 582 418 730 423
rect 582 417 665 418
rect 690 417 730 418
rect 931 406 950 413
rect 983 409 987 542
rect 1126 541 1136 542
rect 1126 537 1178 541
rect 1071 451 1082 466
rect 195 -19 531 -8
rect 515 -40 531 -19
rect 666 -20 673 51
rect 744 -8 758 37
rect 1071 -8 1082 434
rect 1126 423 1136 537
rect 1495 457 1501 546
rect 1331 450 1501 457
rect 1331 448 1338 450
rect 1126 418 1224 423
rect 1126 417 1213 418
rect 1531 413 1535 553
rect 1676 540 1685 553
rect 1676 536 1727 540
rect 1619 447 1633 460
rect 1479 406 1498 413
rect 744 -19 1082 -8
rect 1214 -19 1221 63
rect 1292 -8 1304 37
rect 1619 -8 1633 434
rect 1676 423 1685 536
rect 2042 457 2049 545
rect 1882 451 2049 457
rect 1882 444 1888 451
rect 1676 417 1764 423
rect 1820 407 1830 414
rect 2028 406 2047 413
rect 1292 -19 1633 -8
rect 1765 -18 1772 57
rect 1843 -17 1851 37
rect 1071 -38 1082 -19
rect 1619 -38 1633 -19
<< m2contact >>
rect 55 608 64 615
rect 159 602 165 610
rect 63 553 74 561
rect 600 608 609 615
rect 713 602 722 610
rect 318 528 325 533
rect 167 511 174 519
rect 55 499 61 504
rect 271 503 277 508
rect 299 482 306 489
rect 210 461 221 469
rect 607 553 619 561
rect 1149 603 1158 611
rect 1262 598 1271 606
rect 1809 597 1818 605
rect 234 442 244 449
rect 234 409 244 416
rect 863 528 871 533
rect 712 511 721 526
rect 816 503 825 509
rect 602 498 609 503
rect 844 482 851 489
rect 761 461 770 469
rect 1155 549 1166 558
rect 783 441 790 447
rect 549 406 556 413
rect 783 407 790 414
rect 1412 524 1420 529
rect 1261 507 1270 515
rect 1363 499 1373 505
rect 1149 494 1158 499
rect 1393 473 1400 481
rect 1309 455 1319 465
rect 1331 441 1338 448
rect 1097 407 1104 413
rect 1331 407 1338 414
rect 1703 549 1715 557
rect 1959 523 1968 528
rect 1808 506 1817 514
rect 1911 498 1919 503
rect 1696 493 1704 498
rect 1860 455 1869 464
rect 1882 437 1888 444
rect 1648 406 1655 413
rect 1882 407 1888 414
<< metal2 >>
rect 55 626 174 631
rect 55 615 64 626
rect 159 598 163 602
rect 40 553 63 561
rect 40 425 51 553
rect 158 544 163 598
rect 170 565 174 626
rect 600 625 667 632
rect 600 615 609 625
rect 125 539 163 544
rect 55 534 133 539
rect 55 504 61 534
rect 167 519 174 565
rect 658 563 667 625
rect 1149 622 1205 628
rect 1149 611 1158 622
rect 589 553 607 561
rect 318 507 325 528
rect 277 503 325 507
rect 306 482 556 489
rect 210 425 221 461
rect 40 420 221 425
rect 40 419 115 420
rect 140 419 221 420
rect 210 397 221 419
rect 234 416 244 442
rect 549 413 556 482
rect 589 423 598 553
rect 1696 620 1754 627
rect 713 543 722 602
rect 1696 603 1705 620
rect 602 537 722 543
rect 1132 549 1155 558
rect 602 503 609 537
rect 667 518 712 526
rect 863 507 871 528
rect 825 503 871 507
rect 602 434 609 498
rect 851 482 1104 489
rect 761 423 770 461
rect 589 418 770 423
rect 589 417 665 418
rect 690 417 770 418
rect 761 395 770 417
rect 783 414 790 441
rect 1097 413 1104 482
rect 1132 423 1142 549
rect 1262 540 1271 598
rect 1149 534 1271 540
rect 1679 549 1703 557
rect 1149 499 1158 534
rect 1215 499 1270 507
rect 1412 503 1420 524
rect 1373 499 1420 503
rect 1149 434 1158 494
rect 1400 473 1655 481
rect 1309 423 1319 455
rect 1132 418 1319 423
rect 1132 417 1213 418
rect 1238 417 1319 418
rect 1309 395 1319 417
rect 1331 414 1338 441
rect 1648 413 1655 473
rect 1679 423 1687 549
rect 1809 540 1818 597
rect 1696 532 1818 540
rect 1696 498 1704 532
rect 1763 498 1817 506
rect 1959 502 1968 523
rect 1919 498 1968 502
rect 1696 434 1704 493
rect 1860 423 1869 455
rect 1679 418 1869 423
rect 1679 417 1764 418
rect 1789 417 1869 418
rect 1860 395 1869 417
rect 1882 414 1888 437
<< m3contact >>
rect 1205 622 1215 628
rect 658 549 667 563
rect 1754 620 1763 627
rect 658 518 667 526
rect 602 429 609 434
rect 1205 499 1215 507
rect 1149 429 1158 434
rect 1754 498 1763 506
rect 1696 429 1704 434
<< m123contact >>
rect 193 429 202 434
<< metal3 >>
rect 658 526 667 549
rect 1205 507 1215 622
rect 1754 506 1763 620
rect 202 429 602 434
rect 609 429 1149 434
rect 1158 429 1696 434
use Full_Adder_t2  Full_Adder_t2_0
timestamp 1698872434
transform 0 1 337 -1 0 300
box -125 -337 300 101
use Full_Adder_t2  Full_Adder_t2_1
timestamp 1698872434
transform 0 1 886 -1 0 298
box -125 -337 300 101
use Full_Adder_t2  Full_Adder_t2_2
timestamp 1698872434
transform 0 1 1434 -1 0 298
box -125 -337 300 101
use Full_Adder_t2  Full_Adder_t2_3
timestamp 1698872434
transform 0 1 1985 -1 0 298
box -125 -337 300 101
use XOR  XOR_0 /home/vsoham
timestamp 1698822538
transform 1 0 199 0 1 551
box -144 -89 205 89
use XOR  XOR_1
timestamp 1698822538
transform 1 0 744 0 1 551
box -144 -89 205 89
use XOR  XOR_2
timestamp 1698822538
transform 1 0 1293 0 1 547
box -144 -89 205 89
use XOR  XOR_3
timestamp 1698822538
transform 1 0 1840 0 1 546
box -144 -89 205 89
<< labels >>
flabel metal1 117 -19 124 -7 0 FreeSans 9 0 0 0 S0
flabel metal1 666 -20 673 -6 0 FreeSans 9 0 0 0 S1
flabel metal1 1214 -19 1221 -7 0 FreeSans 9 0 0 0 S2
flabel metal1 1765 -18 1772 -6 0 FreeSans 9 0 0 0 S3
flabel metal1 1843 -17 1851 -5 0 FreeSans 9 0 0 0 C_over
flabel metal1 55 590 64 615 0 FreeSans 9 0 0 0 B0
flabel metal1 600 590 609 615 0 FreeSans 9 0 0 0 B1
flabel metal1 1149 586 1158 611 0 FreeSans 9 0 0 0 B2
flabel metal1 1696 585 1705 610 0 FreeSans 9 0 0 0 B3
flabel metal1 2028 406 2047 413 0 FreeSans 9 0 0 0 A3
flabel metal1 1479 406 1498 413 0 FreeSans 9 0 0 0 A2
flabel metal1 931 406 950 413 0 FreeSans 9 0 0 0 A1
flabel metal1 384 408 403 415 0 FreeSans 9 0 0 0 A0
flabel metal1 17 419 33 425 0 FreeSans 9 0 0 0 VDD
flabel metal1 0 408 7 425 0 FreeSans 9 0 0 0 GND
flabel metal1 163 441 167 445 0 FreeSans 9 0 0 0 C_in
flabel metal1 515 -40 531 -5 0 FreeSans 9 0 0 0 D0
flabel space 1071 -39 1082 -1 0 FreeSans 9 0 0 0 D1
flabel space 1618 -39 1633 -3 0 FreeSans 9 0 0 0 D2
flabel metal1 1071 451 1082 466 0 FreeSans 9 0 0 0 D1
flabel metal1 1619 447 1633 460 0 FreeSans 9 0 0 0 D2
<< end >>
