magic
tech scmos
timestamp 1700128855
<< polysilicon >>
rect 331 -385 409 -378
rect 407 -476 417 -441
<< polycontact >>
rect 319 -385 331 -378
rect 409 -385 419 -378
rect 407 -441 417 -433
rect 407 -484 417 -476
<< metal1 >>
rect 1 168 5 173
rect 350 172 428 181
rect -73 165 5 168
rect 422 164 428 172
rect 729 163 826 166
rect 505 159 609 163
rect 729 159 733 163
rect -106 127 -99 152
rect 758 153 770 158
rect 822 155 826 163
rect -106 123 -90 127
rect -106 109 -99 123
rect -48 111 -41 138
rect 422 117 428 147
rect 822 134 834 139
rect 15 92 20 97
rect -60 89 -53 92
rect -47 89 20 92
rect 379 87 401 90
rect -61 80 -12 83
rect -106 42 -99 49
rect -106 38 -90 42
rect -106 32 -99 38
rect -47 33 -40 53
rect 9 37 13 41
rect -47 26 -32 33
rect -40 25 -32 26
rect -61 4 -53 7
rect -47 4 -12 7
rect -10 4 14 7
rect -64 -6 -15 -3
rect -11 -6 6 -3
rect 1 -15 6 -6
rect -106 -44 -99 -29
rect -106 -48 -90 -44
rect -106 -54 -99 -48
rect -47 -66 -40 -33
rect 396 -53 401 87
rect 408 72 427 77
rect 408 4 414 72
rect 505 62 616 65
rect 408 -15 414 -2
rect 505 -18 589 -14
rect 736 -54 742 -50
rect 453 -71 456 -60
rect -61 -82 -53 -79
rect -47 -82 14 -79
rect 11 -88 14 -82
rect -67 -91 -18 -88
rect -16 -91 -15 -88
rect 11 -91 33 -88
rect 386 -98 421 -95
rect -107 -129 -100 -114
rect -107 -133 -97 -129
rect -107 -140 -100 -133
rect -47 -156 -40 -118
rect -21 -133 -18 -128
rect 53 -130 60 -103
rect 459 -110 463 -89
rect 505 -91 509 -73
rect 663 -72 669 -68
rect 830 -70 834 134
rect 822 -75 834 -70
rect 725 -83 758 -79
rect 505 -95 574 -91
rect 459 -118 493 -110
rect 383 -132 450 -129
rect -64 -167 -53 -164
rect -47 -167 -15 -164
rect 488 -196 504 -193
rect 515 -206 522 -173
rect 538 -183 544 -95
rect 708 -146 715 -124
rect 781 -137 787 -95
rect 820 -142 824 -91
rect 820 -153 836 -142
rect 705 -175 727 -171
rect 538 -187 607 -183
rect 258 -232 263 -223
rect 427 -227 443 -221
rect 258 -237 340 -232
rect 395 -278 400 -228
rect 705 -238 712 -216
rect 722 -263 727 -175
rect 702 -267 756 -263
rect 385 -281 571 -278
rect 53 -303 60 -286
rect 422 -293 428 -281
rect 505 -292 589 -288
rect 752 -307 756 -267
rect 820 -272 824 -153
rect 820 -293 832 -289
rect 229 -361 235 -315
rect 319 -378 331 -341
rect -116 -441 -107 -420
rect 394 -446 402 -329
rect 764 -332 769 -328
rect 614 -364 622 -342
rect 505 -378 611 -375
rect 419 -385 428 -378
rect 407 -430 425 -425
rect 407 -433 417 -430
rect 394 -462 402 -455
rect 505 -458 613 -454
rect 382 -465 402 -462
rect 394 -468 402 -465
rect 394 -473 425 -468
rect 229 -549 235 -497
rect 376 -499 442 -495
rect 827 -497 832 -293
rect 820 -500 832 -497
rect 453 -534 456 -517
rect 237 -549 439 -545
rect 459 -552 463 -538
rect 562 -545 578 -535
rect 752 -534 756 -511
rect 731 -538 756 -534
rect 733 -545 739 -538
rect 480 -549 739 -545
rect 459 -555 747 -552
<< m2contact >>
rect 341 172 350 181
rect -84 162 -78 168
rect 0 152 6 158
rect 422 147 428 152
rect 749 150 758 158
rect -61 121 -54 129
rect 385 129 390 134
rect -12 121 -5 129
rect 504 129 509 134
rect 733 117 740 125
rect -48 105 -41 111
rect 590 93 595 100
rect 766 95 772 101
rect -53 86 -47 92
rect -84 80 -78 86
rect -106 49 -99 57
rect -61 36 -54 44
rect -106 24 -99 32
rect -11 36 -4 44
rect -40 19 -32 25
rect 0 15 6 22
rect -53 1 -47 7
rect -84 -6 -78 0
rect 0 -33 6 -27
rect -61 -50 -54 -42
rect -106 -62 -99 -54
rect -11 -50 -4 -42
rect 699 78 706 83
rect 764 37 771 43
rect 422 27 428 32
rect 734 29 741 36
rect 587 18 592 23
rect 661 14 668 19
rect 408 -2 414 4
rect 699 -3 706 3
rect 408 -21 414 -15
rect 421 -17 428 -11
rect 765 -20 771 -13
rect 442 -41 447 -36
rect -40 -66 -33 -58
rect 301 -61 306 -56
rect 396 -58 401 -53
rect 742 -54 749 -47
rect 453 -60 459 -55
rect 450 -77 456 -71
rect 525 -72 530 -67
rect 570 -72 576 -67
rect 663 -68 669 -63
rect 699 -64 706 -57
rect -53 -85 -47 -79
rect -84 -91 -78 -85
rect 421 -100 428 -95
rect -61 -135 -54 -127
rect -107 -147 -100 -140
rect -27 -133 -21 -128
rect -11 -135 -4 -127
rect 614 -77 623 -68
rect 493 -118 502 -110
rect 53 -137 60 -130
rect 450 -132 456 -126
rect 301 -144 306 -139
rect -40 -156 -30 -148
rect -53 -167 -47 -161
rect 229 -184 235 -178
rect 53 -198 60 -191
rect 483 -196 488 -191
rect 465 -207 470 -202
rect 610 -129 617 -121
rect 781 -144 787 -137
rect 558 -161 567 -154
rect 0 -217 6 -210
rect 610 -221 618 -213
rect 305 -227 310 -221
rect 395 -228 402 -222
rect 421 -227 427 -221
rect 558 -253 567 -246
rect 571 -283 576 -278
rect 53 -309 60 -303
rect 762 -274 771 -266
rect 229 -315 235 -309
rect 0 -353 6 -346
rect 394 -329 402 -321
rect 737 -328 743 -322
rect 764 -328 769 -323
rect 229 -367 235 -361
rect 53 -382 60 -376
rect 0 -398 6 -391
rect 384 -423 389 -418
rect -116 -451 -107 -441
rect 421 -340 428 -335
rect 698 -338 705 -331
rect 524 -346 529 -341
rect 570 -346 575 -341
rect 661 -346 668 -339
rect 614 -372 622 -364
rect 763 -390 769 -384
rect 734 -411 742 -403
rect 504 -423 509 -418
rect 588 -422 593 -417
rect 622 -422 631 -416
rect 661 -430 669 -421
rect 698 -443 705 -437
rect 394 -455 402 -446
rect 762 -447 770 -439
rect 407 -492 417 -484
rect 643 -492 648 -484
rect 229 -497 235 -492
rect 0 -537 6 -529
rect 442 -499 447 -494
rect 733 -500 741 -490
rect 453 -517 459 -512
rect 592 -524 597 -517
rect 439 -549 446 -544
rect 473 -549 480 -544
rect 698 -538 705 -532
rect 779 -549 792 -542
rect 747 -555 756 -549
<< metal2 >>
rect 225 172 341 181
rect -116 -140 -110 162
rect -106 158 -99 172
rect -84 86 -78 162
rect -65 152 0 158
rect 392 147 422 152
rect -61 129 -54 134
rect -61 117 -54 121
rect -12 129 -5 134
rect 390 129 504 134
rect -41 105 -35 111
rect -12 109 -5 121
rect 590 100 595 154
rect 740 117 772 125
rect 766 101 772 117
rect -106 57 -99 66
rect -106 2 -99 24
rect -84 0 -78 80
rect -61 44 -54 49
rect -61 32 -54 36
rect -50 7 -47 86
rect -106 -80 -99 -62
rect -84 -85 -78 -6
rect -61 -42 -54 -37
rect -61 -54 -54 -50
rect -50 -79 -47 1
rect -40 -15 -32 19
rect -61 -127 -54 -122
rect -61 -139 -54 -135
rect -116 -147 -107 -140
rect -107 -391 -100 -147
rect -50 -161 -47 -85
rect -40 -113 -33 -66
rect -27 -128 -24 83
rect -11 44 -4 57
rect -11 11 -4 36
rect 422 23 428 27
rect 6 15 14 22
rect 356 18 587 23
rect -11 6 152 11
rect 0 -27 6 -6
rect 146 0 152 6
rect 269 -7 382 0
rect 414 -2 509 4
rect -11 -42 -4 -29
rect 274 -45 380 -37
rect -11 -54 -4 -50
rect -11 -127 -4 -114
rect 0 -120 146 -112
rect -11 -147 -4 -135
rect -40 -173 -30 -156
rect -66 -181 -30 -173
rect 53 -191 60 -137
rect 301 -139 306 -61
rect 338 -58 396 -53
rect -4 -217 0 -210
rect -33 -353 0 -346
rect 53 -376 60 -309
rect 229 -309 235 -184
rect 338 -221 343 -58
rect 310 -227 343 -221
rect 408 -222 414 -21
rect 349 -321 356 -227
rect 402 -228 414 -222
rect 421 -95 428 -17
rect 447 -41 456 -38
rect 453 -55 456 -41
rect 526 -67 530 18
rect 570 -67 576 -2
rect 661 -7 668 14
rect 699 3 706 78
rect 734 37 764 43
rect 734 36 741 37
rect 618 -22 625 -15
rect 618 -27 669 -22
rect 614 -68 623 -45
rect 663 -63 669 -27
rect 699 -57 706 -3
rect 742 -20 765 -13
rect 742 -47 749 -20
rect 450 -83 456 -77
rect 699 -83 706 -64
rect 450 -88 706 -83
rect 421 -221 427 -100
rect 450 -120 456 -88
rect 502 -117 740 -110
rect 502 -118 606 -117
rect 621 -118 740 -117
rect 450 -126 468 -120
rect 465 -193 468 -126
rect 610 -138 617 -129
rect 610 -144 781 -138
rect 465 -196 483 -193
rect 465 -202 468 -196
rect 349 -329 394 -321
rect 421 -335 427 -227
rect 558 -232 567 -161
rect 610 -204 792 -196
rect 610 -213 618 -204
rect 558 -246 567 -237
rect 756 -274 762 -266
rect 505 -350 512 -323
rect 571 -341 575 -283
rect 626 -323 668 -314
rect 256 -358 512 -350
rect 661 -339 668 -323
rect 743 -328 764 -323
rect -107 -398 0 -391
rect -116 -462 -107 -451
rect 229 -492 235 -367
rect 246 -365 493 -364
rect 255 -373 493 -365
rect 389 -423 504 -418
rect 524 -446 529 -346
rect 578 -373 614 -364
rect 661 -421 669 -398
rect 588 -446 593 -422
rect 402 -455 593 -446
rect 698 -437 705 -338
rect 734 -390 763 -384
rect 734 -403 742 -390
rect 636 -492 643 -484
rect 407 -508 417 -492
rect 447 -498 456 -495
rect 453 -512 456 -498
rect 574 -524 592 -517
rect -66 -537 0 -529
rect 698 -532 705 -443
rect 733 -447 762 -439
rect 733 -490 741 -447
rect 446 -549 473 -545
rect 747 -549 756 -524
rect 784 -542 792 -204
<< m3contact >>
rect -106 172 -99 181
rect 216 172 225 181
rect -116 162 -110 168
rect -72 152 -65 158
rect 590 154 595 159
rect 383 147 392 152
rect -61 134 -54 142
rect -61 109 -54 117
rect -35 105 -29 111
rect 740 150 749 158
rect -106 66 -99 72
rect -61 49 -54 57
rect -61 24 -54 32
rect -61 -37 -54 -29
rect -61 -62 -54 -54
rect -40 -22 -32 -15
rect -61 -122 -54 -114
rect -61 -147 -54 -139
rect -40 -118 -33 -113
rect 14 15 23 22
rect 349 18 356 23
rect 146 -7 152 0
rect 263 -7 269 0
rect 382 -7 388 0
rect 509 -2 515 4
rect 266 -45 274 -37
rect 380 -45 388 -37
rect 0 -108 6 -102
rect 146 -120 155 -112
rect -77 -181 -66 -173
rect -12 -217 -4 -210
rect -40 -353 -33 -346
rect 570 -2 576 4
rect 618 -15 625 -10
rect 661 -15 668 -7
rect 614 -45 623 -37
rect 740 -118 749 -110
rect 558 -237 567 -232
rect 747 -274 756 -266
rect 505 -323 512 -314
rect 618 -323 626 -314
rect 248 -358 256 -350
rect -116 -471 -107 -462
rect 246 -373 255 -365
rect 493 -373 501 -364
rect 570 -373 578 -364
rect 661 -398 669 -389
rect 622 -416 631 -406
rect 407 -517 417 -508
rect -77 -537 -66 -529
rect 747 -524 756 -517
<< m123contact >>
rect -106 152 -99 158
rect 641 125 646 133
rect 625 18 630 23
rect 349 -227 356 -221
rect 340 -237 345 -232
rect 319 -341 331 -333
<< metal3 >>
rect -99 172 216 181
rect -110 163 405 168
rect 398 159 405 163
rect -99 152 -72 158
rect 398 155 590 159
rect -89 134 -61 142
rect 15 135 646 142
rect 641 133 646 135
rect -97 109 -61 117
rect -29 105 0 111
rect -99 66 -44 72
rect -97 49 -61 57
rect -89 24 -61 32
rect -8 12 0 105
rect 283 30 630 38
rect 14 12 23 15
rect -8 6 23 12
rect -32 -22 6 -15
rect -97 -37 -61 -29
rect -97 -62 -61 -54
rect -61 -98 -54 -62
rect -97 -122 -61 -114
rect -97 -147 -61 -139
rect -116 -545 -107 -471
rect -97 -517 -89 -147
rect -77 -484 -66 -181
rect -40 -333 -33 -118
rect -12 -186 -4 -88
rect 0 -102 6 -22
rect 14 -171 23 6
rect 152 -7 263 0
rect 249 -45 266 -37
rect 155 -120 211 -112
rect 202 -153 211 -120
rect 202 -160 216 -153
rect 283 -186 293 30
rect 625 23 630 30
rect 315 4 331 14
rect -12 -192 293 -186
rect -12 -210 -4 -192
rect 319 -333 331 4
rect 349 -221 356 18
rect 388 -7 494 0
rect 515 -2 570 4
rect 487 -10 494 -7
rect 487 -15 618 -10
rect 650 -15 661 -7
rect 388 -45 614 -37
rect 740 -110 749 150
rect 345 -237 558 -232
rect 539 -263 549 -237
rect 512 -323 618 -314
rect -77 -529 -66 -492
rect -55 -541 -48 -345
rect -40 -341 278 -333
rect -40 -346 -33 -341
rect 226 -358 248 -350
rect 271 -389 278 -341
rect 501 -373 570 -364
rect 271 -398 661 -389
rect 560 -416 622 -406
rect 747 -517 756 -274
rect 407 -541 417 -517
rect -55 -548 417 -541
<< m234contact >>
rect -12 134 -5 142
rect -27 83 -22 88
rect -106 -6 -99 2
rect 0 -6 6 2
rect -11 -62 -4 -54
rect -106 -88 -99 -80
rect 628 -492 636 -484
rect 567 -524 574 -517
<< m4contact >>
rect 376 147 383 152
rect -97 134 -89 142
rect 8 135 15 142
rect -44 66 -38 72
rect -97 24 -89 32
rect -61 -105 -54 -98
rect -12 -88 -4 -80
rect -97 -524 -89 -517
rect 241 -45 249 -37
rect 216 -160 226 -153
rect 14 -178 23 -171
rect 303 4 315 14
rect 642 -15 650 -7
rect 539 -275 549 -263
rect -77 -492 -66 -484
rect -55 -345 -48 -338
rect -116 -555 -107 -545
rect 216 -358 226 -350
rect 238 -373 246 -365
rect 551 -416 560 -406
<< metal4 >>
rect -97 158 -43 164
rect -12 163 383 171
rect -97 142 -89 158
rect -12 142 -5 163
rect 16 148 315 155
rect 8 88 15 135
rect -22 83 15 88
rect -38 66 211 72
rect 203 36 211 66
rect 203 29 249 36
rect -97 15 -89 24
rect -116 7 -89 15
rect -116 -365 -110 7
rect -99 -6 0 2
rect 241 -37 249 29
rect 303 14 315 148
rect 376 152 383 163
rect 258 -15 642 -7
rect 258 -54 266 -15
rect -4 -62 266 -54
rect -99 -88 -12 -80
rect -54 -105 265 -98
rect -55 -178 14 -171
rect -55 -338 -48 -178
rect 216 -350 226 -160
rect -116 -373 238 -365
rect 257 -406 265 -105
rect 539 -391 549 -275
rect 257 -416 551 -406
rect -66 -492 628 -484
rect -89 -524 567 -517
rect -107 -555 539 -545
<< m5contact >>
rect -43 158 -38 164
rect 10 148 16 155
rect 539 -400 549 -391
rect 539 -555 549 -545
<< metal5 >>
rect -38 158 16 164
rect 10 155 16 158
rect 539 -545 549 -400
use XNOR  XNOR_3
timestamp 1699700809
transform 1 0 291 0 1 -519
box -291 -33 98 145
use XNOR  XNOR_2
timestamp 1699700809
transform 1 0 291 0 1 -335
box -291 -33 98 145
use 4_input  4_input_1
timestamp 1699636190
transform 1 0 604 0 1 -330
box 0 0 1 1
use 3in_AND  3in_AND_1
timestamp 1698787690
transform 1 0 643 0 1 -407
box 0 0 1 1
use AND_2  AND_2_1
timestamp 1698776759
transform 1 0 598 0 1 -501
box -8 -37 143 47
use 5_input_AND  5_input_AND_1
timestamp 1699638001
transform 0 1 467 -1 0 -292
box -12 -45 256 42
use 4_input_OR  4_input_OR_1
timestamp 1699703636
transform 0 1 788 -1 0 -271
box 226 32 235 36
use XNOR  XNOR_1
timestamp 1699700809
transform 1 0 291 0 1 -152
box -291 -33 98 145
use 5_input_AND  5_input_AND_2
timestamp 1699638001
transform 1 0 262 0 1 -182
box -12 -45 256 42
use CMOS_in  CMOS_in_5
timestamp 1699269643
transform 1 0 -34 0 1 -42
box -13 -40 30 39
use CMOS_in  CMOS_in_4
timestamp 1699269643
transform 1 0 -84 0 1 -42
box -13 -40 30 39
use CMOS_in  CMOS_in_6
timestamp 1699269643
transform 1 0 -84 0 1 -127
box -13 -40 30 39
use CMOS_in  CMOS_in_7
timestamp 1699269643
transform 1 0 -34 0 1 -127
box -13 -40 30 39
use XNOR  XNOR_0
timestamp 1699700809
transform 1 0 291 0 1 33
box -291 -33 98 145
use CMOS_in  CMOS_in_3
timestamp 1699269643
transform 1 0 -34 0 1 44
box -13 -40 30 39
use CMOS_in  CMOS_in_2
timestamp 1699269643
transform 1 0 -84 0 1 44
box -13 -40 30 39
use 4_input  4_input_0
timestamp 1699636190
transform 1 0 605 0 1 -56
box 0 0 1 1
use AND_2  AND_2_3
timestamp 1698776759
transform 1 0 568 0 1 -230
box -8 -37 143 47
use AND_2  AND_2_2
timestamp 1698776759
transform 1 0 568 0 1 -138
box -8 -37 143 47
use 5_input_AND  5_input_AND_0
timestamp 1699638001
transform 0 1 467 -1 0 165
box -12 -45 256 42
use 4_input_OR  4_input_OR_0
timestamp 1699703636
transform 0 1 790 -1 0 156
box 226 32 235 36
use CMOS_in  CMOS_in_1
timestamp 1699269643
transform 1 0 -35 0 1 129
box -13 -40 30 39
use CMOS_in  CMOS_in_0
timestamp 1699269643
transform 1 0 -84 0 1 129
box -13 -40 30 39
use 3in_AND  3in_AND_0
timestamp 1698787690
transform 1 0 642 0 1 33
box 0 0 1 1
use AND_2  AND_2_0
timestamp 1698776759
transform 1 0 596 0 1 116
box -8 -37 143 47
<< labels >>
flabel metal1 -106 123 -99 127 0 FreeSans 9 0 0 0 A0
flabel metal1 -48 123 -41 127 0 FreeSans 9 0 0 0 B0
flabel metal1 -106 38 -99 42 0 FreeSans 9 0 0 0 A1
flabel metal1 -47 38 -40 42 0 FreeSans 9 0 0 0 B1
flabel metal1 -106 -48 -99 -44 0 FreeSans 9 0 0 0 A2
flabel metal1 -47 -48 -40 -44 0 FreeSans 9 0 0 0 B2
flabel metal1 -107 -133 -100 -129 0 FreeSans 9 0 0 0 A3
flabel metal1 -47 -133 -40 -129 0 FreeSans 9 0 0 0 B3
flabel metal1 -116 -436 -107 -420 0 FreeSans 9 0 0 0 En
flabel metal1 820 -153 836 -142 0 FreeSans 9 0 0 0 VDD
flabel metal1 562 -549 578 -535 0 FreeSans 9 0 0 0 GND
flabel metal1 708 -133 715 -124 0 FreeSans 9 0 0 0 Gth
flabel metal1 705 -224 712 -216 0 FreeSans 9 0 0 0 Lth
flabel metal1 515 -190 522 -186 0 FreeSans 9 0 0 0 Eql
<< end >>
