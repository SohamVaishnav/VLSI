magic
tech scmos
timestamp 1699703636
<< labels >>
flabel metal1 226 32 235 36 0 FreeSans 9 0 0 0 VDD
<< end >>
