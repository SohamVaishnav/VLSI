magic
tech scmos
timestamp 1698778229
<< metal1 >>
rect -80 84 -77 89
rect 61 85 85 89
rect -135 81 -120 84
rect -96 81 -77 84
rect -31 51 -24 59
rect 68 43 77 47
rect -144 39 -129 43
rect -97 39 -84 42
rect -89 26 -84 39
rect -89 19 -73 26
rect -129 5 -121 8
rect -99 5 -94 8
rect -5 5 0 9
rect -99 2 0 5
rect -81 -7 -75 -2
rect -135 -10 -119 -7
rect -96 -10 -75 -7
rect 73 -18 77 43
rect 82 32 85 85
rect 194 -4 205 -1
rect 73 -23 87 -18
rect 119 -23 125 -18
rect -32 -40 -25 -32
rect 65 -48 78 -44
rect -144 -52 -129 -48
rect -101 -52 -84 -49
rect -89 -65 -84 -52
rect -89 -72 -74 -65
rect 100 -82 104 -30
rect -130 -86 -118 -83
rect -97 -86 -94 -83
rect -6 -86 -1 -82
rect 63 -86 104 -82
rect -97 -89 -1 -86
use OR_2  OR_2_0 /home/vsoham
timestamp 1698776833
transform 1 0 129 0 1 -2
box -47 -31 71 40
use AND_2  AND_2_1 /home/vsoham
timestamp 1698776759
transform 1 0 -73 0 1 -49
box -8 -37 143 47
use AND_2  AND_2_0
timestamp 1698776759
transform 1 0 -72 0 1 42
box -8 -37 143 47
use CMOS_in  CMOS_in_1 /home/vsoham
timestamp 1698776633
transform 1 0 -124 0 1 -46
box -13 -40 30 39
use CMOS_in  CMOS_in_0
timestamp 1698776633
transform 1 0 -124 0 1 45
box -13 -40 30 39
<< labels >>
flabel metal1 -144 -52 -137 -48 0 FreeSans 9 0 0 0 B
flabel metal1 -144 39 -137 43 0 FreeSans 9 0 0 0 A
flabel metal1 194 -4 205 -1 0 FreeSans 9 0 0 0 OUT
flabel metal1 65 -48 78 -44 0 FreeSans 9 0 0 0 ABc
flabel metal1 119 -23 125 -18 0 FreeSans 9 0 0 0 ABc
flabel metal1 -31 51 -24 59 0 FreeSans 9 0 0 0 B
flabel metal1 -32 -40 -25 -32 0 FreeSans 9 0 0 0 A
flabel metal1 -135 81 -123 84 0 FreeSans 9 0 0 0 VDD
flabel metal1 -135 -10 -123 -7 0 FreeSans 9 0 0 0 VDD
flabel metal1 -130 -86 -118 -83 0 FreeSans 9 0 0 0 GND
flabel metal1 -129 5 -121 8 0 FreeSans 9 0 0 0 GND
<< end >>
