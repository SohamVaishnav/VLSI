magic
tech scmos
timestamp 1700523696
<< polysilicon >>
rect 1385 639 1393 652
rect 1385 635 2120 639
rect 2114 607 2120 635
<< polycontact >>
rect 1385 652 1393 658
rect 2114 601 2120 607
<< metal1 >>
rect 887 856 893 865
rect 1486 855 1513 861
rect 1486 844 1492 855
rect 1569 844 1592 850
rect 19 820 25 829
rect 466 820 472 829
rect 1573 804 1580 808
rect 2223 786 2241 793
rect 1670 741 1676 745
rect 1737 741 1743 745
rect 1804 741 1810 745
rect 1871 741 1877 745
rect 1670 705 1676 709
rect 1737 705 1743 709
rect 1804 705 1810 709
rect 1860 705 1866 709
rect 1931 662 1935 674
rect 2019 666 2023 674
rect 2107 666 2111 674
rect 2195 666 2199 674
rect 1294 645 1302 658
rect 887 615 893 624
rect 1207 619 1300 622
rect 1318 619 1322 648
rect 1638 627 1643 646
rect 1726 642 1743 646
rect 1790 642 1807 646
rect 1863 642 1873 646
rect 1882 628 1886 653
rect 2157 645 2163 646
rect 2157 638 2179 645
rect 2237 629 2241 653
rect 1207 605 1210 619
rect 1266 565 1271 572
rect 2114 571 2120 601
rect 2212 599 2220 606
rect 2212 515 2220 522
rect 1266 481 1271 488
rect 2212 415 2220 422
rect 1260 388 1271 393
rect 887 377 893 386
rect 1260 381 1266 388
rect 19 365 25 374
rect 467 365 473 374
rect 2212 325 2220 332
rect 2171 315 2183 321
rect 1260 304 1271 309
rect 1262 297 1266 304
rect 1892 191 1904 197
rect 887 132 893 141
rect 1892 107 1904 113
rect 1220 7 1224 59
rect 1220 3 1536 7
<< m2contact >>
rect 1939 735 1947 746
rect 2027 735 2037 744
rect 2115 735 2123 742
rect 2203 735 2211 742
rect 1970 686 1977 693
rect 2058 686 2065 693
rect 2146 686 2153 693
rect 2234 686 2241 693
rect 1893 646 1899 652
rect 1981 646 1987 652
rect 2069 646 2075 652
rect 2157 646 2163 652
<< metal2 >>
rect 1345 869 1904 877
rect 1244 855 1498 861
rect 1244 774 1252 855
rect 1492 844 1498 855
rect 1895 833 1904 869
rect 1895 824 2211 833
rect 1220 764 1252 774
rect 1336 703 1345 791
rect 1939 746 1947 810
rect 2027 744 2037 810
rect 2115 742 2123 800
rect 2203 742 2211 824
rect 1199 696 1345 703
rect 1199 688 1208 696
rect 861 681 1208 688
rect 1977 686 2058 693
rect 2065 686 2146 693
rect 2153 686 2234 693
rect 1518 668 1648 677
rect 1662 609 1670 677
rect 1819 668 1922 677
rect 1916 652 1922 668
rect 1899 646 1981 652
rect 1987 646 2069 652
rect 2075 646 2157 652
rect 1641 602 1670 609
rect 1641 506 1651 602
rect 1622 495 1651 506
rect 864 194 1208 201
rect 424 16 433 145
rect 424 8 671 16
<< m3contact >>
rect 1939 810 1948 819
rect 2027 810 2037 819
rect 1210 764 1220 774
rect 854 681 861 688
rect 854 194 864 201
rect 1208 194 1217 201
rect 671 8 679 16
<< m123contact >>
rect 1573 797 1580 804
rect 1907 786 1914 793
rect 1665 777 1672 786
rect 1995 786 2002 793
rect 2083 786 2090 793
rect 2171 786 2178 793
rect 1294 638 1302 645
rect 366 591 373 600
rect 813 593 820 600
rect 366 137 374 145
rect 814 138 821 147
<< metal3 >>
rect 431 887 1642 895
rect 431 600 440 887
rect 1631 819 1642 887
rect 2027 819 2037 828
rect 1631 810 1939 819
rect 1580 797 1914 804
rect 1907 793 1914 797
rect 1914 786 1995 793
rect 2002 786 2083 793
rect 2090 786 2171 793
rect 1643 780 1665 786
rect 1306 777 1665 780
rect 1306 773 1651 777
rect 1210 718 1219 764
rect 871 711 1219 718
rect 854 600 861 681
rect 373 591 440 600
rect 820 593 861 600
rect 1208 201 1217 665
rect 1306 645 1314 773
rect 1302 638 1314 645
rect 854 147 864 194
rect 374 137 433 145
rect 821 138 864 147
rect 671 38 1231 45
rect 671 16 679 38
<< m234contact >>
rect 1336 869 1345 877
rect 1336 791 1345 799
rect 2115 800 2123 808
<< m4contact >>
rect 1208 665 1217 672
<< metal4 >>
rect 1242 893 1391 900
rect 1242 770 1251 893
rect 1384 884 1391 893
rect 1384 877 1703 884
rect 1336 799 1345 869
rect 1694 847 1703 877
rect 1694 837 1983 847
rect 1976 808 1983 837
rect 1976 800 2115 808
rect 1208 762 1251 770
rect 1208 672 1217 762
<< m345contact >>
rect 2027 828 2037 836
rect 1231 38 1242 47
<< metal5 >>
rect 1231 873 1679 882
rect 1231 47 1242 873
rect 1668 836 1679 873
rect 1668 828 2027 836
use 4_bit_ANDer_t2  4_bit_ANDer_t2_0
timestamp 1700522344
transform 0 1 1822 -1 0 781
box -5 -201 139 64
use 4_bit_Adder_t3  4_bit_Adder_t3_0
timestamp 1700521624
transform 1 0 290 0 1 554
box -290 -554 950 348
use 4_bit_Comp_t2  4_bit_Comp_t2_0
timestamp 1700522019
transform 1 0 1375 0 1 464
box -122 -463 895 168
use Decoder  Decoder_0
timestamp 1700521764
transform 0 1 1440 -1 0 692
box -158 -188 50 169
use AND_2  AND_2_3
timestamp 1698776759
transform 0 1 2194 -1 0 785
box -8 -37 143 47
use AND_2  AND_2_2
timestamp 1698776759
transform 0 1 2106 -1 0 785
box -8 -37 143 47
use AND_2  AND_2_1
timestamp 1698776759
transform 0 1 2018 -1 0 785
box -8 -37 143 47
use AND_2  AND_2_0
timestamp 1698776759
transform 0 1 1930 -1 0 785
box -8 -37 143 47
<< labels >>
flabel metal1 1931 666 1935 674 0 FreeSans 9 0 0 0 S3
flabel metal1 2019 666 2023 674 0 FreeSans 9 0 0 0 S2
flabel metal1 2107 666 2111 674 0 FreeSans 9 0 0 0 S1
flabel metal1 2195 666 2199 674 0 FreeSans 9 0 0 0 S0
flabel metal1 1498 855 1513 861 0 FreeSans 9 0 0 0 Sel1
flabel metal1 1577 844 1592 850 0 FreeSans 9 0 0 0 Sel0
flabel metal1 1863 642 1873 646 0 FreeSans 9 0 0 0 C0
flabel metal1 1797 642 1807 646 0 FreeSans 9 0 0 0 C1
flabel metal1 1733 642 1743 646 0 FreeSans 9 0 0 0 C2
flabel metal1 1638 627 1643 635 0 FreeSans 9 0 0 0 C3
flabel metal1 2223 786 2237 793 0 FreeSans 9 0 0 0 VDD
flabel metal1 2157 638 2179 645 0 FreeSans 9 0 0 0 GND
flabel metal1 2171 315 2183 321 0 FreeSans 9 0 0 0 Eql
flabel metal1 1892 191 1904 197 0 FreeSans 9 0 0 0 Lth
flabel metal1 1892 107 1904 113 0 FreeSans 9 0 0 0 Gth
flabel metal1 1266 565 1271 572 0 FreeSans 9 0 0 0 A3
flabel metal1 1266 481 1271 488 0 FreeSans 9 0 0 0 B3
flabel metal1 1260 381 1266 388 0 FreeSans 9 0 0 0 A2
flabel metal1 1262 297 1266 304 0 FreeSans 9 0 0 0 B2
flabel metal1 2212 599 2220 606 0 FreeSans 9 0 0 0 A0
flabel metal1 2212 515 2220 522 0 FreeSans 9 0 0 0 B0
flabel metal1 2212 415 2220 422 0 FreeSans 9 0 0 0 A1
flabel metal1 2212 325 2220 332 0 FreeSans 9 0 0 0 B1
flabel metal1 1804 705 1810 709 0 FreeSans 9 0 0 0 B1
flabel metal1 1804 741 1810 745 0 FreeSans 9 0 0 0 A1
flabel metal1 1871 741 1877 745 0 FreeSans 9 0 0 0 A0
flabel metal1 1860 705 1866 709 0 FreeSans 9 0 0 0 B0
flabel metal1 1737 741 1743 745 0 FreeSans 9 0 0 0 A2
flabel metal1 1737 705 1743 709 0 FreeSans 9 0 0 0 B2
flabel metal1 1670 741 1676 745 0 FreeSans 9 0 0 0 A3
flabel metal1 1670 705 1676 709 0 FreeSans 9 0 0 0 B3
flabel metal1 887 856 893 865 0 FreeSans 9 0 0 0 B0
flabel metal1 887 615 893 624 0 FreeSans 9 0 0 0 B1
flabel metal1 887 377 893 386 0 FreeSans 9 0 0 0 B2
flabel metal1 887 132 893 141 0 FreeSans 9 0 0 0 B3
flabel metal1 19 820 25 829 0 FreeSans 9 0 0 0 A3
flabel metal1 19 365 25 374 0 FreeSans 9 0 0 0 A2
flabel metal1 467 365 473 374 0 FreeSans 9 0 0 0 A1
flabel metal1 466 820 472 829 0 FreeSans 9 0 0 0 A0
<< end >>
