magic
tech scmos
timestamp 1700515345
use Decoder  Decoder_0
timestamp 1699864537
transform 0 1 1440 -1 0 692
box -158 -188 50 169
use 4_bit_Comp_t2  4_bit_Comp_t2_0
timestamp 1700501889
transform 1 0 1375 0 1 464
box -122 -463 895 168
use 4_bit_Adder_t3  4_bit_Adder_t3_0
timestamp 1699914285
transform 1 0 290 0 1 554
box -290 -554 950 348
<< end >>
