magic
tech scmos
timestamp 1698711931
<< nwell >>
rect -1 -4 28 38
rect 42 -4 71 38
rect 86 -4 115 38
rect 130 -4 159 38
rect 174 -4 203 38
rect 219 -4 248 38
<< ntransistor >>
rect 12 -29 14 -17
rect 55 -29 57 -17
rect 99 -29 101 -17
rect 143 -29 145 -17
rect 187 -29 189 -17
rect 232 -29 234 -17
<< ptransistor >>
rect 6 14 20 18
rect 49 14 63 18
rect 93 14 107 18
rect 137 14 151 18
rect 181 14 195 18
rect 226 14 240 18
<< ndiffusion >>
rect 10 -29 12 -17
rect 14 -29 16 -17
rect 53 -29 55 -17
rect 57 -29 59 -17
rect 97 -29 99 -17
rect 101 -29 103 -17
rect 141 -29 143 -17
rect 145 -29 147 -17
rect 185 -29 187 -17
rect 189 -29 191 -17
rect 230 -29 232 -17
rect 234 -29 236 -17
<< pdiffusion >>
rect 6 18 20 21
rect 49 18 63 21
rect 93 18 107 21
rect 137 18 151 21
rect 181 18 195 21
rect 226 18 240 21
rect 6 12 20 14
rect 49 12 63 14
rect 93 12 107 14
rect 137 12 151 14
rect 181 12 195 14
rect 226 12 240 14
<< ndcontact >>
rect 4 -29 10 -17
rect 16 -29 22 -17
rect 47 -29 53 -17
rect 59 -29 65 -17
rect 91 -29 97 -17
rect 103 -29 109 -17
rect 135 -29 141 -17
rect 147 -29 153 -17
rect 179 -29 185 -17
rect 191 -29 197 -17
rect 224 -29 230 -17
rect 236 -29 242 -17
<< pdcontact >>
rect 6 21 20 30
rect 49 21 63 30
rect 93 21 107 30
rect 137 21 151 30
rect 181 21 195 30
rect 226 21 240 30
rect 6 3 20 12
rect 49 3 63 12
rect 93 3 107 12
rect 137 3 151 12
rect 181 3 195 12
rect 226 3 240 12
<< polysilicon >>
rect -12 14 6 18
rect 20 14 28 18
rect 35 14 49 18
rect 63 14 71 18
rect 80 14 93 18
rect 107 14 115 18
rect 125 14 137 18
rect 151 14 159 18
rect 168 14 181 18
rect 195 14 203 18
rect 213 14 226 18
rect 240 14 248 18
rect -12 -32 -8 14
rect 12 -17 14 -14
rect 12 -32 14 -29
rect 35 -32 39 14
rect 55 -17 57 -14
rect 55 -32 57 -29
rect 80 -32 84 14
rect 99 -17 101 -14
rect 99 -32 101 -29
rect 125 -32 129 14
rect 143 -17 145 -14
rect 143 -32 145 -29
rect 168 -32 172 14
rect 213 -3 217 14
rect 187 -17 189 -14
rect 187 -32 189 -29
rect 213 -32 217 -9
rect 232 -17 234 -14
rect 232 -32 234 -29
rect -12 -35 -4 -32
rect 1 -35 15 -32
rect 35 -35 43 -32
rect 48 -35 58 -32
rect 80 -35 88 -32
rect 93 -35 102 -32
rect 125 -35 133 -32
rect 138 -35 146 -32
rect 168 -35 176 -32
rect 181 -35 190 -32
rect 213 -35 235 -32
<< polycontact >>
rect 211 -9 217 -3
rect -4 -39 1 -32
rect 43 -39 48 -32
rect 88 -39 93 -32
rect 133 -39 138 -32
rect 176 -39 181 -32
<< metal1 >>
rect -6 38 248 42
rect 11 30 15 38
rect 54 30 58 38
rect 98 30 102 38
rect 142 30 146 38
rect 186 30 190 38
rect 231 30 235 38
rect 11 -4 15 3
rect 54 -4 58 3
rect 98 -4 102 3
rect 142 -4 146 3
rect 186 -4 190 3
rect -5 -8 211 -4
rect -5 -21 -1 -8
rect 231 -4 235 3
rect 231 -8 256 -4
rect 237 -14 242 -11
rect 237 -17 240 -14
rect -5 -25 4 -21
rect 22 -25 47 -21
rect 65 -25 91 -21
rect 109 -25 135 -21
rect 153 -25 179 -21
rect 197 -25 206 -21
rect 203 -30 206 -25
rect -4 -45 1 -39
rect 43 -45 48 -39
rect 88 -45 93 -39
rect 133 -45 138 -39
rect 176 -45 181 -39
rect 226 -39 229 -29
rect 245 -39 248 -8
rect 226 -45 248 -39
<< labels >>
flabel metal1 -2 38 202 42 0 FreeSans 8 0 0 0 VDD
flabel metal1 176 -45 181 -41 0 FreeSans 9 0 0 0 E
flabel metal1 133 -45 138 -41 0 FreeSans 9 0 0 0 D
flabel metal1 88 -45 93 -41 0 FreeSans 9 0 0 0 C
flabel metal1 43 -45 48 -41 0 FreeSans 9 0 0 0 B
flabel metal1 -4 -45 1 -41 0 FreeSans 9 0 0 0 A
flabel metal1 237 -14 242 -11 0 FreeSans 8 0 0 0 GND
flabel metal1 248 -8 256 -4 0 FreeSans 8 0 0 0 OUT
flabel metal1 197 -25 206 -21 0 FreeSans 8 0 0 0 GND
<< end >>
