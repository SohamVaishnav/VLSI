magic
tech scmos
timestamp 1700132798
<< nwell >>
rect -45 -10 -19 25
rect -9 -10 17 25
rect 27 -10 53 25
rect 64 -10 90 25
<< ntransistor >>
rect -38 -28 -26 -23
rect -2 -28 10 -23
rect 34 -28 46 -23
rect 71 -28 83 -23
<< ptransistor >>
rect -38 6 -26 10
rect -2 6 10 10
rect 34 6 46 10
rect 71 6 83 10
<< ndiffusion >>
rect -38 -23 -26 -22
rect -2 -23 10 -22
rect 34 -23 46 -22
rect 71 -23 83 -22
rect -38 -29 -26 -28
rect -2 -29 10 -28
rect 34 -29 46 -28
rect 71 -29 83 -28
<< pdiffusion >>
rect -38 10 -26 11
rect -2 10 10 11
rect 34 10 46 11
rect 71 10 83 11
rect -38 4 -26 6
rect -2 4 10 6
rect 34 4 46 6
rect 71 4 83 6
<< ndcontact >>
rect -38 -22 -26 -16
rect -2 -22 10 -16
rect 34 -22 46 -16
rect 71 -22 83 -16
rect -38 -35 -26 -29
rect -2 -35 10 -29
rect 34 -35 46 -29
rect 71 -35 83 -29
<< pdcontact >>
rect -38 11 -26 18
rect -2 11 10 18
rect 34 11 46 18
rect 71 11 83 18
rect -38 -3 -26 4
rect -2 -3 10 4
rect 34 -3 46 4
rect 71 -3 83 4
<< polysilicon >>
rect -41 6 -38 10
rect -26 6 -19 10
rect -45 -23 -41 5
rect -5 6 -2 10
rect 10 6 17 10
rect -9 -23 -5 5
rect 31 6 34 10
rect 46 6 53 10
rect 64 6 71 10
rect 83 6 90 10
rect 27 -23 31 5
rect 64 -6 68 6
rect 64 -23 68 -10
rect -45 -28 -38 -23
rect -26 -28 -19 -23
rect -9 -28 -2 -23
rect 10 -28 17 -23
rect 27 -28 34 -23
rect 46 -28 53 -23
rect 64 -28 71 -23
rect 83 -28 90 -23
<< polycontact >>
rect -45 5 -41 10
rect -9 5 -5 10
rect 27 5 31 10
rect 64 -10 68 -6
<< metal1 >>
rect -45 21 90 25
rect -34 18 -30 21
rect 2 18 6 21
rect 38 18 42 21
rect 75 18 79 21
rect -49 5 -45 10
rect -13 5 -9 10
rect 23 5 27 10
rect -34 -6 -30 -3
rect 2 -6 6 -3
rect 38 -6 42 -3
rect 75 -6 79 -3
rect 86 -6 90 2
rect -34 -10 64 -6
rect 75 -10 90 -6
rect -34 -16 -30 -10
rect 75 -16 79 -10
rect 10 -21 34 -17
rect 86 -17 90 -10
rect -34 -39 6 -35
rect 38 -39 90 -35
<< end >>
