magic
tech scmos
timestamp 1698872434
<< metal1 >>
rect -125 97 141 101
rect -125 -34 -119 97
rect -102 54 -96 97
rect 115 58 118 97
rect -115 -7 -108 49
rect 267 17 293 21
rect 214 8 243 11
rect -97 -22 -85 -19
rect 231 -31 281 -28
rect -125 -37 -87 -34
rect -125 -129 -119 -37
rect -116 -103 -109 -49
rect 212 -60 293 -57
rect 83 -75 108 -69
rect -97 -113 -84 -110
rect -125 -132 -87 -129
rect -125 -220 -119 -132
rect 261 -142 270 -120
rect -116 -201 -109 -144
rect 258 -152 293 -149
rect -97 -208 -92 -205
rect 217 -220 252 -213
rect -125 -223 -86 -220
rect -125 -232 -119 -223
rect -114 -230 -92 -226
rect -114 -261 -109 -230
rect 223 -246 293 -243
rect 80 -261 102 -256
rect -109 -265 -104 -261
rect -97 -299 -86 -296
rect -104 -330 -97 -299
rect -115 -333 -97 -330
rect 214 -333 293 -329
rect -115 -337 293 -333
<< m2contact >>
rect 178 63 183 71
rect 252 55 257 60
rect 2 24 11 32
rect 127 31 132 38
rect -103 12 -96 17
rect 293 12 300 21
rect 243 4 250 11
rect -115 -15 -108 -7
rect -104 -25 -97 -19
rect 281 -35 289 -28
rect -116 -49 -109 -42
rect 152 -50 161 -45
rect 1 -67 10 -59
rect 293 -66 300 -57
rect 108 -75 117 -69
rect -104 -113 -97 -107
rect 147 -142 152 -137
rect 188 -142 193 -137
rect 1 -162 10 -154
rect 293 -158 300 -149
rect -116 -208 -109 -201
rect -104 -208 -97 -202
rect -92 -231 -87 -226
rect 151 -236 160 -231
rect 0 -253 9 -245
rect 293 -252 300 -243
rect 102 -261 110 -256
rect 266 -261 271 -256
rect -114 -270 -109 -261
rect 192 -287 197 -279
rect -104 -299 -97 -293
rect 266 -295 271 -290
rect 141 -319 146 -312
rect 293 -337 300 -329
<< metal2 >>
rect -103 91 132 97
rect -103 17 -96 91
rect 2 32 11 76
rect 127 38 132 91
rect 178 71 183 91
rect 225 55 252 59
rect -108 -15 -84 -7
rect -116 -42 -109 -26
rect -104 -107 -97 -25
rect -93 -30 -84 -15
rect 2 -19 11 24
rect -93 -37 10 -30
rect 1 -59 10 -37
rect 152 -69 161 -50
rect 117 -75 161 -69
rect 225 -87 231 55
rect 243 -77 250 4
rect -116 -211 -109 -208
rect -104 -202 -97 -113
rect 188 -93 231 -87
rect 188 -137 193 -93
rect 147 -154 152 -142
rect 147 -160 263 -154
rect 1 -199 10 -162
rect -10 -203 10 -199
rect -10 -206 -4 -203
rect -114 -312 -109 -270
rect -104 -293 -97 -208
rect -57 -210 -4 -206
rect -57 -226 -49 -210
rect -87 -230 -49 -226
rect 0 -245 9 -217
rect 0 -261 9 -253
rect 102 -221 160 -215
rect 102 -256 110 -221
rect 151 -231 160 -221
rect 256 -222 263 -160
rect 241 -227 263 -222
rect 241 -228 247 -227
rect 281 -246 289 -35
rect 141 -249 289 -246
rect 293 -57 300 12
rect 293 -149 300 -66
rect 293 -243 300 -158
rect 0 -268 98 -261
rect 89 -299 98 -268
rect 141 -312 146 -249
rect 192 -295 197 -287
rect 241 -290 247 -268
rect 241 -295 266 -290
rect -114 -319 141 -312
rect 293 -329 300 -252
<< m3contact >>
rect 2 76 11 84
rect 178 91 183 97
rect -116 -26 -109 -19
rect 2 -26 11 -19
rect -116 -217 -109 -211
rect 0 -217 9 -211
rect 241 -233 247 -228
rect 89 -306 98 -299
rect 271 -261 279 -256
rect 241 -268 247 -263
rect 192 -302 197 -295
<< m123contact >>
rect 243 -84 250 -77
<< metal3 >>
rect 2 91 178 97
rect 2 84 11 91
rect -109 -26 2 -19
rect 250 -84 279 -77
rect -109 -217 0 -211
rect 241 -263 247 -233
rect 271 -256 279 -84
rect 110 -299 192 -295
rect 98 -302 192 -299
rect 98 -306 110 -302
use XOR  XOR_0 /home/vsoham
timestamp 1698822538
transform 1 0 33 0 1 -27
box -144 -89 205 89
use XOR  XOR_1
timestamp 1698822538
transform 1 0 32 0 1 -213
box -144 -89 205 89
use OR_2  OR_2_0 /home/vsoham
timestamp 1698776833
transform 1 0 194 0 1 -121
box -47 -31 71 40
use AND_2  AND_2_0 /home/vsoham
timestamp 1698776759
transform 1 0 133 0 1 54
box -8 -37 143 47
use AND_2  AND_2_1
timestamp 1698776759
transform 1 0 147 0 1 -296
box -8 -37 143 47
<< end >>
