magic
tech scmos
timestamp 1698858438
<< metal1 >>
rect -11 85 -4 93
rect -239 50 -233 53
rect 148 51 161 70
rect -239 47 -224 50
rect 129 47 164 51
rect -247 9 -245 10
rect -247 5 -236 9
rect -223 -29 -222 -24
rect 91 -38 96 -22
rect -239 -44 -231 -39
rect 109 -64 118 13
rect 86 -67 118 -64
rect 130 -75 174 -71
rect -257 -82 -256 -77
rect -34 -82 -25 -77
rect -257 -86 -235 -82
rect 136 -113 158 -108
rect -225 -120 -224 -115
rect -228 -138 -227 -132
rect -265 -223 -257 -148
rect 86 -156 87 -151
rect -245 -177 -241 -172
rect 171 -175 174 -75
rect 91 -220 101 -217
rect -265 -226 -231 -223
rect 92 -229 101 -220
rect 81 -249 109 -246
rect -243 -264 -234 -263
rect -37 -264 -28 -259
rect -256 -268 -234 -264
rect -23 -277 -19 -250
rect 79 -292 85 -260
rect 135 -292 138 -283
rect -240 -302 -215 -299
rect -33 -303 -28 -294
rect -17 -303 -12 -294
rect 79 -296 138 -292
<< m2contact >>
rect 42 55 47 66
rect 164 41 173 51
rect -9 23 -4 30
rect -232 -29 -223 -24
rect 96 -38 102 -32
rect 5 -75 12 -70
rect -265 -86 -257 -77
rect -232 -120 -225 -115
rect -28 -120 -17 -114
rect -3 -120 3 -115
rect 148 -122 158 -113
rect -239 -138 -228 -132
rect 80 -156 86 -151
rect -135 -165 -126 -157
rect 116 -175 125 -165
rect -43 -215 -34 -206
rect 116 -212 121 -207
rect -136 -256 -127 -248
rect -23 -250 -18 -245
rect -23 -282 -18 -277
rect -28 -303 -17 -294
<< metal2 >>
rect -21 97 47 102
rect -21 72 -16 97
rect -265 66 -134 72
rect -125 66 -16 72
rect 42 66 47 97
rect -265 -77 -257 66
rect -253 58 -4 62
rect -253 10 -247 58
rect -9 30 -4 58
rect -234 -26 -232 -24
rect -253 -29 -232 -26
rect -253 -117 -249 -29
rect -21 -71 -16 -47
rect 96 -68 102 -38
rect -21 -75 5 -71
rect 58 -75 102 -68
rect 58 -101 63 -75
rect -233 -117 -232 -115
rect -253 -120 -232 -117
rect -239 -142 -228 -138
rect -257 -148 -228 -142
rect -135 -172 -126 -165
rect -241 -213 -233 -177
rect -188 -177 -126 -172
rect -188 -203 -181 -177
rect -28 -206 -17 -120
rect -3 -151 1 -120
rect -3 -155 80 -151
rect 79 -156 80 -155
rect 148 -152 158 -122
rect 94 -160 158 -152
rect -241 -221 -127 -213
rect -34 -215 -17 -206
rect -136 -248 -127 -221
rect -28 -245 -17 -215
rect -28 -250 -23 -245
rect -18 -250 -17 -245
rect 12 -234 20 -169
rect 94 -209 104 -160
rect 164 -165 173 41
rect 125 -175 173 -165
rect 114 -209 116 -207
rect 94 -212 116 -209
rect 12 -239 15 -234
rect -181 -264 -179 -263
rect 12 -264 20 -239
rect -181 -268 20 -264
rect -28 -282 -23 -278
rect -18 -282 -17 -278
rect -28 -294 -17 -282
<< m3contact >>
rect -11 85 -4 93
rect -134 66 -125 72
rect -239 47 -233 53
rect -134 17 -125 25
rect -239 -44 -233 -39
rect -25 -47 -16 -41
rect -135 -74 -126 -66
rect 16 -57 25 -52
rect -34 -82 -25 -77
rect -188 -209 -181 -203
rect 7 -141 12 -134
rect 12 -169 20 -163
rect 15 -239 24 -234
rect -241 -268 -234 -263
rect -188 -268 -181 -263
rect -33 -264 -26 -259
<< m123contact >>
rect -253 5 -247 10
rect 58 -109 63 -101
rect -265 -148 -257 -142
rect -241 -177 -233 -172
<< metal3 >>
rect -11 80 -4 85
rect -239 76 -4 80
rect -239 53 -233 76
rect -265 47 -239 53
rect -265 -142 -257 47
rect -253 -126 -247 5
rect -239 -39 -233 47
rect -134 25 -125 66
rect -21 -41 -16 76
rect 16 -64 25 -57
rect -135 -126 -126 -74
rect -34 -67 25 -64
rect -34 -77 -25 -67
rect -253 -134 -126 -126
rect 7 -169 12 -141
rect -233 -173 -229 -172
rect 58 -173 63 -109
rect -233 -177 63 -173
rect -188 -263 -181 -209
rect -234 -264 -232 -263
rect -190 -264 -188 -263
rect -234 -268 -188 -264
rect 15 -260 24 -239
rect -26 -264 24 -260
use OR_2  OR_2_0
timestamp 1698776833
transform 0 1 137 -1 0 -217
box -47 -31 71 40
use XOR  XOR_1
timestamp 1698822538
transform 1 0 -104 0 1 -216
box -144 -89 205 89
use AND_2  AND_2_1
timestamp 1698776759
transform 1 0 13 0 1 -118
box -8 -37 143 47
use AND_2  AND_2_0
timestamp 1698776759
transform 1 0 -3 0 1 46
box -8 -37 143 47
use XOR  XOR_0
timestamp 1698822538
transform 1 0 -103 0 1 -34
box -144 -89 205 89
<< labels >>
flabel metal1 -247 5 -241 9 0 FreeSans 9 0 0 0 A
flabel metal1 -247 -86 -241 -82 0 FreeSans 9 0 0 0 B
flabel metal1 79 -270 85 -260 0 FreeSans 9 0 0 0 Carry
flabel metal1 -256 -268 -248 -264 0 FreeSans 9 0 0 0 C
flabel metal1 -240 -302 -230 -299 0 FreeSans 9 0 0 0 GND
flabel metal1 -265 -165 -257 -148 0 FreeSans 9 0 0 0 VDD
flabel metal1 148 47 161 70 0 FreeSans 9 0 0 0 AB
flabel metal1 91 -32 96 -22 0 FreeSans 9 0 0 0 AxB
flabel metal1 136 -113 158 -108 0 FreeSans 9 0 0 0 C(AxB)
flabel metal1 92 -229 101 -217 0 FreeSans 9 0 0 0 Sum
<< end >>
