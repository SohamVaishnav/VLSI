magic
tech scmos
timestamp 1698959774
<< polysilicon >>
rect -671 245 -660 631
rect -208 245 -198 633
rect 249 245 261 631
rect 708 246 720 632
rect -671 236 -651 245
rect -208 236 -189 245
rect 249 236 270 245
rect 708 236 729 246
<< polycontact >>
rect -671 631 -660 642
rect -208 633 -198 643
rect 249 631 261 640
rect 708 632 720 641
rect -651 236 -644 245
rect -189 236 -182 245
rect 270 236 277 245
rect 729 236 736 246
<< metal1 >>
rect 484 657 492 667
rect 944 657 952 667
rect -671 648 -401 656
rect -208 649 67 657
rect 249 649 495 657
rect 708 649 955 657
rect -671 642 -660 648
rect -660 583 -653 622
rect -420 609 -414 648
rect -208 643 -198 649
rect -420 603 -317 609
rect -353 591 -261 594
rect -660 492 -653 522
rect -274 440 -261 591
rect -198 583 -191 623
rect 42 610 54 649
rect 249 640 261 649
rect 708 641 720 649
rect 118 591 201 594
rect -223 561 -172 564
rect -223 529 -214 561
rect -223 473 -214 523
rect -198 492 -191 524
rect -223 470 -167 473
rect 188 440 201 591
rect 261 583 268 623
rect 582 591 660 594
rect 248 561 289 564
rect 248 473 255 561
rect 261 494 268 526
rect 248 470 293 473
rect 649 440 660 591
rect 720 582 727 622
rect 1033 591 1118 594
rect 699 561 754 564
rect 699 473 705 561
rect 720 492 727 525
rect 699 470 756 473
rect -274 436 -180 440
rect 188 436 287 440
rect 646 436 738 440
rect 1108 436 1118 591
rect -650 388 -643 396
rect -188 381 -181 396
rect 271 388 278 396
rect 730 388 737 396
rect -591 314 -583 320
rect -129 314 -120 320
rect 330 314 337 320
rect 789 314 798 320
rect -224 210 -214 226
rect 234 214 244 230
rect -274 202 -214 210
rect 188 206 244 214
rect 691 213 701 229
rect 647 205 701 213
rect 1115 197 1129 204
rect -671 169 -664 174
rect -289 119 -269 126
rect 179 119 193 126
rect 638 119 652 126
rect 1097 119 1111 126
rect -660 94 -654 110
rect -658 2 -647 9
rect -242 2 -173 9
rect 220 2 289 9
rect 679 2 748 9
<< m2contact >>
rect 495 649 507 657
rect 955 649 964 657
rect -445 640 -439 645
rect -547 607 -538 615
rect 16 640 23 645
rect -317 603 -310 609
rect -660 576 -653 583
rect -455 550 -449 556
rect -317 552 -310 561
rect -397 533 -388 538
rect -660 522 -653 530
rect -548 516 -539 524
rect -325 523 -318 529
rect -449 508 -438 514
rect -660 484 -653 492
rect -591 461 -583 470
rect -85 607 -76 615
rect 475 640 482 645
rect 937 640 943 645
rect 42 602 54 610
rect -198 577 -191 583
rect 6 550 13 556
rect 145 552 152 561
rect 65 533 74 538
rect -223 523 -214 529
rect -198 524 -191 531
rect -86 516 -77 524
rect 13 508 24 513
rect -198 485 -191 492
rect -129 460 -120 470
rect 374 607 383 615
rect 261 577 268 583
rect 465 550 472 556
rect 604 552 612 562
rect 524 533 533 538
rect 261 526 268 532
rect 373 516 382 524
rect 472 508 483 514
rect 261 486 268 494
rect 330 461 337 470
rect 833 607 842 615
rect 720 576 727 582
rect 925 550 931 556
rect 1063 552 1071 562
rect 983 533 992 538
rect 720 525 727 531
rect 832 516 841 524
rect 931 508 942 514
rect 720 485 727 492
rect 789 462 798 470
rect -591 320 -583 327
rect -129 320 -120 326
rect 330 320 337 326
rect 789 320 798 326
rect -214 202 -204 210
rect 244 206 255 214
rect 701 205 712 213
rect -651 188 -644 195
rect -189 176 -182 185
rect 270 183 277 192
rect 729 185 736 195
rect -671 164 -664 169
rect -651 165 -644 170
<< metal2 >>
rect -660 560 -653 576
rect -660 555 -551 560
rect -660 530 -653 543
rect -558 524 -551 555
rect -547 550 -538 607
rect -445 556 -439 640
rect -449 550 -439 556
rect -317 561 -310 603
rect -198 560 -191 577
rect -198 553 -89 560
rect -558 516 -548 524
rect -397 514 -388 533
rect -198 531 -191 543
rect -318 523 -223 529
rect -96 524 -89 553
rect -85 549 -76 607
rect 16 556 23 640
rect 54 602 152 610
rect 13 550 23 556
rect 145 561 152 602
rect 261 561 268 577
rect 261 555 370 561
rect -96 516 -86 524
rect -438 508 -388 514
rect 65 513 74 533
rect 261 532 268 543
rect 363 524 370 555
rect 374 549 383 607
rect 475 556 482 640
rect 495 607 507 649
rect 495 598 612 607
rect 472 550 482 556
rect 604 562 612 598
rect 720 561 727 576
rect 720 554 829 561
rect 363 516 373 524
rect 524 514 533 533
rect 720 531 727 543
rect 822 524 829 554
rect 833 549 842 607
rect 937 556 943 640
rect 955 607 964 649
rect 955 598 1071 607
rect 931 550 943 556
rect 1063 562 1071 598
rect 822 516 832 524
rect 983 514 992 533
rect 24 508 74 513
rect 483 508 533 514
rect 942 508 992 514
rect -660 461 -653 484
rect -660 447 -653 454
rect -671 440 -653 447
rect -591 449 -583 461
rect -198 461 -191 485
rect -129 451 -120 460
rect 261 461 268 486
rect 330 447 337 461
rect 720 461 727 485
rect 789 455 798 462
rect -671 195 -660 440
rect -591 327 -583 415
rect -129 326 -120 415
rect 330 326 337 415
rect 789 326 798 414
rect -671 188 -651 195
rect -214 185 -204 202
rect 244 192 255 206
rect 701 195 712 205
rect -214 176 -189 185
rect 244 183 270 192
rect 701 185 729 195
rect -664 165 -651 169
<< m3contact >>
rect -660 543 -653 550
rect -547 543 -538 550
rect -198 543 -191 549
rect -85 543 -76 549
rect 261 543 268 549
rect 374 543 383 549
rect 720 543 727 549
rect 833 543 842 549
rect -660 454 -653 461
rect -198 454 -191 461
rect -591 443 -583 449
rect 261 454 268 461
rect -129 443 -120 451
rect 720 454 727 461
rect 789 447 798 455
rect 330 440 337 447
rect -591 415 -583 422
rect -129 415 -120 423
rect 330 415 337 423
rect 789 414 798 423
<< m123contact >>
rect -458 561 -451 569
rect -437 470 -429 480
<< metal3 >>
rect -451 561 -429 569
rect -653 543 -547 550
rect -437 480 -429 561
rect -191 543 -85 549
rect 268 543 374 549
rect 727 543 833 549
rect -653 454 -198 461
rect -191 455 261 461
rect -191 454 -133 455
rect -116 454 261 455
rect 268 454 720 461
rect -591 422 -583 443
rect -129 423 -120 443
rect 330 423 337 440
rect 789 423 798 447
use XOR  XOR_3 /home/vsoham
timestamp 1698822538
transform 1 0 -516 0 1 556
box -144 -89 205 89
use XOR  XOR_2
timestamp 1698822538
transform 1 0 -54 0 1 556
box -144 -89 205 89
use XOR  XOR_1
timestamp 1698822538
transform 1 0 405 0 1 556
box -144 -89 205 89
use XOR  XOR_0
timestamp 1698822538
transform 1 0 864 0 1 556
box -144 -89 205 89
use Full_Adder_t2  Full_Adder_t2_3
timestamp 1698872434
transform 1 0 845 0 1 339
box -125 -337 300 101
use Full_Adder_t2  Full_Adder_t2_2
timestamp 1698872434
transform 1 0 386 0 1 339
box -125 -337 300 101
use Full_Adder_t2  Full_Adder_t2_1
timestamp 1698872434
transform 1 0 -73 0 1 339
box -125 -337 300 101
use Full_Adder_t2  Full_Adder_t2_0
timestamp 1698872434
transform 1 0 -535 0 1 339
box -125 -337 300 101
<< labels >>
flabel metal1 -671 169 -664 174 0 FreeSans 9 0 0 0 C_in
flabel metal1 -658 2 -651 9 0 FreeSans 9 0 0 0 GND
flabel metal1 -660 94 -654 106 0 FreeSans 9 0 0 0 VDD
flabel metal1 -188 388 -181 396 0 FreeSans 9 0 0 0 A1
flabel metal1 271 388 278 396 0 FreeSans 9 0 0 0 A2
flabel metal1 730 388 737 396 0 FreeSans 9 0 0 0 A3
flabel metal1 720 614 727 622 0 FreeSans 9 0 0 0 B3
flabel metal1 261 615 268 623 0 FreeSans 9 0 0 0 B2
flabel metal1 -198 615 -191 623 0 FreeSans 9 0 0 0 B1
flabel metal1 -660 614 -653 622 0 FreeSans 9 0 0 0 B0
flabel metal1 -650 388 -643 396 0 FreeSans 9 0 0 0 A0
flabel metal1 -283 119 -269 126 0 FreeSans 9 0 0 0 S0
flabel metal1 179 119 193 126 0 FreeSans 9 0 0 0 S1
flabel metal1 638 119 652 126 0 FreeSans 9 0 0 0 S2
flabel metal1 1097 119 1111 126 0 FreeSans 9 0 0 0 S3
flabel metal1 1115 197 1129 204 0 FreeSans 9 0 0 0 C_over
flabel metal1 -414 648 -401 656 0 FreeSans 9 0 0 0 b_eff0
flabel metal1 54 649 67 657 0 FreeSans 9 0 0 0 b_eff1
flabel metal1 484 649 492 667 0 FreeSans 9 0 0 0 b_eff2
flabel metal1 944 649 952 667 0 FreeSans 9 0 0 0 b_eff3
flabel metal1 -224 210 -214 226 0 FreeSans 9 0 0 0 D0
flabel metal1 234 214 244 230 0 FreeSans 9 0 0 0 D1
flabel metal1 691 213 701 229 0 FreeSans 9 0 0 0 D2
<< end >>
