* SPICE3 file created from Full_Adder_t3.ext - technology: scmos

.option scale=0.09u

M1000 VDD OR_2_0/a_n35_n16# C_out OR_2_0/w_40_n2# pfet w=15 l=5
+  ad=4554 pd=1516 as=135 ps=48
M1001 OR_2_0/a_n35_n16# m1_295_n32# GND Gnd nfet w=15 l=5
+  ad=210 pd=88 as=3609 ps=1252
M1002 OR_2_0/a_n35_n16# m1_295_n32# OR_2_0/a_n35_5# OR_2_0/w_n1_n2# pfet w=15 l=5
+  ad=135 pd=48 as=270 ps=96
M1003 C_out OR_2_0/a_n35_n16# GND Gnd nfet w=15 l=5
+  ad=105 pd=44 as=0 ps=0
M1004 VDD m1_252_n34# OR_2_0/a_n35_5# OR_2_0/w_n42_n2# pfet w=15 l=5
+  ad=0 pd=0 as=0 ps=0
M1005 OR_2_0/a_n35_n16# m1_252_n34# GND Gnd nfet w=15 l=5
+  ad=0 pd=0 as=0 ps=0
M1006 VDD C AND_2_1/a_9_10# AND_2_1/w_n1_1# pfet w=20 l=7
+  ad=0 pd=0 as=360 ps=116
M1007 AND_2_1/a_9_10# C AND_2_1/a_10_n33# Gnd nfet w=18 l=7
+  ad=180 pd=56 as=360 ps=112
M1008 VDD AND_2_1/a_9_10# m1_252_n34# AND_2_1/w_101_1# pfet w=20 l=7
+  ad=0 pd=0 as=180 ps=58
M1009 AND_2_1/a_10_n33# m1_0_n50# GND Gnd nfet w=18 l=7
+  ad=0 pd=0 as=0 ps=0
M1010 VDD m1_0_n50# AND_2_1/a_9_10# AND_2_1/w_50_1# pfet w=20 l=7
+  ad=0 pd=0 as=0 ps=0
M1011 m1_252_n34# AND_2_1/a_9_10# GND Gnd nfet w=18 l=7
+  ad=180 pd=56 as=0 ps=0
M1012 VDD A AND_2_0/a_9_10# AND_2_0/w_n1_1# pfet w=20 l=7
+  ad=0 pd=0 as=360 ps=116
M1013 AND_2_0/a_9_10# A AND_2_0/a_10_n33# Gnd nfet w=18 l=7
+  ad=180 pd=56 as=360 ps=112
M1014 VDD AND_2_0/a_9_10# m1_295_n32# AND_2_0/w_101_1# pfet w=20 l=7
+  ad=0 pd=0 as=180 ps=58
M1015 AND_2_0/a_10_n33# B GND Gnd nfet w=18 l=7
+  ad=0 pd=0 as=0 ps=0
M1016 VDD B AND_2_0/a_9_10# AND_2_0/w_50_1# pfet w=20 l=7
+  ad=0 pd=0 as=0 ps=0
M1017 m1_295_n32# AND_2_0/a_9_10# GND Gnd nfet w=18 l=7
+  ad=180 pd=56 as=0 ps=0
M1018 VDD XOR_0/OR_2_0/a_n35_n16# m1_0_n50# XOR_0/OR_2_0/w_40_n2# pfet w=15 l=5
+  ad=0 pd=0 as=135 ps=48
M1019 XOR_0/OR_2_0/a_n35_n16# XOR_0/m1_65_n48# GND Gnd nfet w=15 l=5
+  ad=210 pd=88 as=0 ps=0
M1020 XOR_0/OR_2_0/a_n35_n16# XOR_0/m1_65_n48# XOR_0/OR_2_0/a_n35_5# XOR_0/OR_2_0/w_n1_n2# pfet w=15 l=5
+  ad=135 pd=48 as=270 ps=96
M1021 m1_0_n50# XOR_0/OR_2_0/a_n35_n16# GND Gnd nfet w=15 l=5
+  ad=105 pd=44 as=0 ps=0
M1022 VDD XOR_0/m1_68_43# XOR_0/OR_2_0/a_n35_5# XOR_0/OR_2_0/w_n42_n2# pfet w=15 l=5
+  ad=0 pd=0 as=0 ps=0
M1023 XOR_0/OR_2_0/a_n35_n16# XOR_0/m1_68_43# GND Gnd nfet w=15 l=5
+  ad=0 pd=0 as=0 ps=0
M1024 XOR_0/m1_n97_39# A GND Gnd nfet w=14 l=4
+  ad=126 pd=46 as=0 ps=0
M1025 VDD A XOR_0/m1_n97_39# XOR_0/CMOS_in_0/w_0_0# pfet w=14 l=4
+  ad=0 pd=0 as=126 ps=46
M1026 VDD XOR_0/m1_n97_39# XOR_0/AND_2_0/a_9_10# XOR_0/AND_2_0/w_n1_1# pfet w=20 l=7
+  ad=0 pd=0 as=360 ps=116
M1027 XOR_0/AND_2_0/a_9_10# XOR_0/m1_n97_39# XOR_0/AND_2_0/a_10_n33# Gnd nfet w=18 l=7
+  ad=180 pd=56 as=360 ps=112
M1028 VDD XOR_0/AND_2_0/a_9_10# XOR_0/m1_68_43# XOR_0/AND_2_0/w_101_1# pfet w=20 l=7
+  ad=0 pd=0 as=180 ps=58
M1029 XOR_0/AND_2_0/a_10_n33# B GND Gnd nfet w=18 l=7
+  ad=0 pd=0 as=0 ps=0
M1030 VDD B XOR_0/AND_2_0/a_9_10# XOR_0/AND_2_0/w_50_1# pfet w=20 l=7
+  ad=0 pd=0 as=0 ps=0
M1031 XOR_0/m1_68_43# XOR_0/AND_2_0/a_9_10# GND Gnd nfet w=18 l=7
+  ad=180 pd=56 as=0 ps=0
M1032 VDD XOR_0/m1_n101_n52# XOR_0/AND_2_1/a_9_10# XOR_0/AND_2_1/w_n1_1# pfet w=20 l=7
+  ad=0 pd=0 as=360 ps=116
M1033 XOR_0/AND_2_1/a_9_10# XOR_0/m1_n101_n52# XOR_0/AND_2_1/a_10_n33# Gnd nfet w=18 l=7
+  ad=180 pd=56 as=360 ps=112
M1034 VDD XOR_0/AND_2_1/a_9_10# XOR_0/m1_65_n48# XOR_0/AND_2_1/w_101_1# pfet w=20 l=7
+  ad=0 pd=0 as=180 ps=58
M1035 XOR_0/AND_2_1/a_10_n33# A GND Gnd nfet w=18 l=7
+  ad=0 pd=0 as=0 ps=0
M1036 VDD A XOR_0/AND_2_1/a_9_10# XOR_0/AND_2_1/w_50_1# pfet w=20 l=7
+  ad=0 pd=0 as=0 ps=0
M1037 XOR_0/m1_65_n48# XOR_0/AND_2_1/a_9_10# GND Gnd nfet w=18 l=7
+  ad=180 pd=56 as=0 ps=0
M1038 XOR_0/m1_n101_n52# B GND Gnd nfet w=14 l=4
+  ad=126 pd=46 as=0 ps=0
M1039 VDD B XOR_0/m1_n101_n52# XOR_0/CMOS_in_1/w_0_0# pfet w=14 l=4
+  ad=0 pd=0 as=126 ps=46
M1040 VDD XOR_1/OR_2_0/a_n35_n16# Sum XOR_1/OR_2_0/w_40_n2# pfet w=15 l=5
+  ad=0 pd=0 as=135 ps=48
M1041 XOR_1/OR_2_0/a_n35_n16# XOR_1/m1_65_n48# GND Gnd nfet w=15 l=5
+  ad=210 pd=88 as=0 ps=0
M1042 XOR_1/OR_2_0/a_n35_n16# XOR_1/m1_65_n48# XOR_1/OR_2_0/a_n35_5# XOR_1/OR_2_0/w_n1_n2# pfet w=15 l=5
+  ad=135 pd=48 as=270 ps=96
M1043 Sum XOR_1/OR_2_0/a_n35_n16# GND Gnd nfet w=15 l=5
+  ad=105 pd=44 as=0 ps=0
M1044 VDD XOR_1/m1_68_43# XOR_1/OR_2_0/a_n35_5# XOR_1/OR_2_0/w_n42_n2# pfet w=15 l=5
+  ad=0 pd=0 as=0 ps=0
M1045 XOR_1/OR_2_0/a_n35_n16# XOR_1/m1_68_43# GND Gnd nfet w=15 l=5
+  ad=0 pd=0 as=0 ps=0
M1046 XOR_1/m1_n97_39# m1_0_n50# GND Gnd nfet w=14 l=4
+  ad=126 pd=46 as=0 ps=0
M1047 VDD m1_0_n50# XOR_1/m1_n97_39# XOR_1/CMOS_in_0/w_0_0# pfet w=14 l=4
+  ad=0 pd=0 as=126 ps=46
M1048 VDD XOR_1/m1_n97_39# XOR_1/AND_2_0/a_9_10# XOR_1/AND_2_0/w_n1_1# pfet w=20 l=7
+  ad=0 pd=0 as=360 ps=116
M1049 XOR_1/AND_2_0/a_9_10# XOR_1/m1_n97_39# XOR_1/AND_2_0/a_10_n33# Gnd nfet w=18 l=7
+  ad=180 pd=56 as=360 ps=112
M1050 VDD XOR_1/AND_2_0/a_9_10# XOR_1/m1_68_43# XOR_1/AND_2_0/w_101_1# pfet w=20 l=7
+  ad=0 pd=0 as=180 ps=58
M1051 XOR_1/AND_2_0/a_10_n33# C GND Gnd nfet w=18 l=7
+  ad=0 pd=0 as=0 ps=0
M1052 VDD C XOR_1/AND_2_0/a_9_10# XOR_1/AND_2_0/w_50_1# pfet w=20 l=7
+  ad=0 pd=0 as=0 ps=0
M1053 XOR_1/m1_68_43# XOR_1/AND_2_0/a_9_10# GND Gnd nfet w=18 l=7
+  ad=180 pd=56 as=0 ps=0
M1054 VDD XOR_1/m1_n101_n52# XOR_1/AND_2_1/a_9_10# XOR_1/AND_2_1/w_n1_1# pfet w=20 l=7
+  ad=0 pd=0 as=360 ps=116
M1055 XOR_1/AND_2_1/a_9_10# XOR_1/m1_n101_n52# XOR_1/AND_2_1/a_10_n33# Gnd nfet w=18 l=7
+  ad=180 pd=56 as=360 ps=112
M1056 VDD XOR_1/AND_2_1/a_9_10# XOR_1/m1_65_n48# XOR_1/AND_2_1/w_101_1# pfet w=20 l=7
+  ad=0 pd=0 as=180 ps=58
M1057 XOR_1/AND_2_1/a_10_n33# m1_0_n50# GND Gnd nfet w=18 l=7
+  ad=0 pd=0 as=0 ps=0
M1058 VDD m1_0_n50# XOR_1/AND_2_1/a_9_10# XOR_1/AND_2_1/w_50_1# pfet w=20 l=7
+  ad=0 pd=0 as=0 ps=0
M1059 XOR_1/m1_65_n48# XOR_1/AND_2_1/a_9_10# GND Gnd nfet w=18 l=7
+  ad=180 pd=56 as=0 ps=0
M1060 XOR_1/m1_n101_n52# C GND Gnd nfet w=14 l=4
+  ad=126 pd=46 as=0 ps=0
M1061 VDD C XOR_1/m1_n101_n52# XOR_1/CMOS_in_1/w_0_0# pfet w=14 l=4
+  ad=0 pd=0 as=126 ps=46
C0 A B 2.21fF
C1 VDD GND 5.62fF
C2 VDD Gnd 3.44fF
C3 C Gnd 3.05fF
C4 m1_0_n50# Gnd 3.47fF
C5 GND Gnd 7.40fF
C6 B Gnd 3.42fF
C7 A Gnd 3.12fF
