magic
tech scmos
timestamp 1698787690
<< end >>
