module Nor_G(Y, A, B);
    input A, B;
    output Y, C;
    Or_G G(C, A, B);
    assign Y = ~C;
endmodule